`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SzDRgzu7qVyBB50Gxp58VQ2J2gsvF9/dbD8XAfcwjoBBEvrcs4ca6znodWInS5XXMXOK+tae5QyR
NC/XIZGbqw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eAdPhBHsXTGh5vzT0lOk8RLFoFi6/bhEzdby9Qk/00aje4YrGXP9CItMf+9Ddy5tjTS6PHmkBbfv
raNlY4NrUxpeSkYHRVnZrudlkD2M0uhKw5CJ9DypalNFsTHNJYic3pS4j58hzDJI0to3SuGdcUDz
v2nAtjvVT0hTBoOBctU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vgz93PAqLHJIk2ulPw0igqbp19viwtBROP4kHq/91uZeaIe6HRetjeu8S3kNpUEC2GzbG8nS4QZo
BbIgLHMqqu91QuhaO7pyVfBgFlKmL5b5rQ3A4/4W8U1O5A3dC4iUkOh4m7m2TcwuYuY4VmzHdOB7
ONDvgHpRpbA8jY/02RITuDMin9DnFYqBBqxQOPFYGpGSqawC2iG4/C07LG4V7q+SyCXSsjkQ5CDZ
W3g8W5KZLsLB+3vZnwy42J8LA/+umE3aHWBFlWiYbwXngfpAvNgpB0GvKZYOsuX4B3x6sH/Yhhc8
z1A5nQjYVQ+9DuplEGIFr/+gkjkOX5p2HhVtCg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tmBQ05yQXHGH3+Gn4eFEjAiU0o5eT7VWgFM4QSmfSMTFuLvsnNAJLkscyGbF7iK2RC1nB02rjuJV
KWPlvG968PcxEsKoCXOp+zeDOzndWx/aQOXcIVx32A/7IsNGL20YGUlcSlwTseOHcttr8jSvJfwk
dKEL5jK9G/WEi8pkvFLGXLH1lCU+RLDp7HeNGY2Lea+Xy+/2XDB5htDyUSXFxhsy0cu3UsEASV00
SXRnW3r1MXcMVwhYnKmH9cVFIfgtj6cRgvRQG4BDzmziCksj/QHzYBmM7G2v0i4kSOJ20+yNMovT
X7I8Q0Kq76S2pbBeeFGCMOnwu/h6UgYd/xib/A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lssvx0lk+DkoCNIS12XWbXhRHt0SHPN+N2dvqJho9DNT1sNN+kpSUobmQUmqVilV9Lh7+z7VBtul
lWg3crXNGO5gotJqO8GUEQoSCjcm5rEzO27J8NbZ0ZE28YZELKnPWd1FF6Uxnx669kwl1dC2j6Tp
S2lo6Aj5/zQ0BQEOAz2jLZvTeTLrQ8HMG5VfKVIRPWzexLnggVDVt5aQXUDwzRprIp4tr0EZOUm4
tWlqYKPheo4Q+oXITR4D3LQBVExLodPWIx5LZmw2c947PrET5gzBJN4c965eUuEpJqY3pw8F2LPT
AbeZ9ePx11JJWFR+u10wo3pAeTaF9Tno2LDO5w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oR+01AVFGS8kZ3pCNoM0CVB4qctAgs1h1qboHJJjJl2DNE5q7GP3bsw0FFi+KRktMYqdhMNeu/ct
DCqPqeKoMj/BAuN8nZ8l1g8n6wH0+opy9UWrhNXvHXVYhulaj4MSpJ8CkVpEwMYol6bWr+MgN6R0
yi8lVDFnue0GCYMiMuM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WRqhaHOwzYTMhqaui33AtC+ejGSAexd4kULR+vSjKepoWb5iul+uAhxy/JPeLgQj7Xu3oXsNDdmP
DDNthRf9IbW7cB7Jz1cRbWwT5BnIjbRGIzFlByrUzB4QCHQO9x3zTkhGVXPPVQThTEeypq8Jqsdo
dzeewNiFhIfKWQGEauEog8jOSuZnvr1q5PMk0Tte1yGjH8arFWfrpe9t25bLajClYt3QzUa+OtBb
2s8u0hPn5OnEo5Cd3+vI++Ytaal5TjMqtgQH9wGZWp6aezag4QKOnTT97sHsFvZZdLhNTq+5zxon
xWDvmAISS6rlyaTLRcTjWVN3pO+qbCdOzITDsg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 63104)
`protect data_block
o0c/crRrYF58CmLEEWAB6mZAFoXostQn9dv8RjgQwoJBg1jEJf1zeSrzYM05Hel0M2PuuFwXUiJB
OWv0tPQvjfROTcF3cG7eG82RHF0Jv058K7N2rqWtWroQ+zogfRvsWfI63V6ielCw2xvwBuJWEveV
eVWXf6Yp5R2OT0hVCz4WVCvsu6qNOD1OMGokNHRIrjiXwOrb748AxdJRxchV3o9ZkoRA9BGv1Qod
Qs5JuvWzq4En85QZnzVIwpsK6HqTfNzEYEtw3xH1n7Wt8POCEo+RB8bpPblQ2xMgPU7lopqU4Mvr
eA1IAq6wJwhT7uDvDkf+HKGCaaWwkhz2wPlq9LaUckdYRFSijOlbS6wqO0yAte+pqyCsJLoJzP7W
TYa2kih9bbPRKYVBpaGL9qk6El29md/EujMqtej/Z7/yXgji4Gw2GPR7BjExaYoGBO+yG7pnNA8B
kE9oJveJVV8g3daBbAaJfa7EhCDyYsJdNv3zre1PAfdvRvW/cLlu6vGbK05CeMAyR2ujsR/KYq5I
cJD/Apj7/LpLVzRCFlsY4DU8NMGMvBGCDDpnFAg5UvT1pQyX7b3tdy5n2lRN34egxaXWjiiwvFIz
DWSVsk3eQTnOEhH7LwfjiSWR03iGRHYQeqCkm6S+A7BArznTryMskC3FN6nL2q7VJIG2GYXUBdcN
zdX81tUBXvdyyXn5inT5fMxZeHSNewrC2p3LwS8Vuzm3e7yIsD7daNMKo8A8q8OqDSOX9ZsERNkC
IB7NQQiFcg9R85gTmtMLWpS70JeFGLW8k0kKeZcUoXVYHQ4gXJNH68Cc7xQGHqt46nehPWuLfMbd
gUqCyfqCOk9YWgFsfxzFbAq3QyKewLYC/Swxk7KZXSEflhF8pd1ypNBmXxkLEd71FMKjaX+gd2l0
3F9eNEAl/xcoOcUVnoX0ceOsnCKPS5LodPsHnk3IaKkmddlqAL3lEWL+TVZhmv9Vaijln6jbCHyk
tF8USc6mmpAjL7KKg/ycAsNJw2jlRbtb/tvLUfclMRZ7Yob1EFh2aaDW/24JK+yYK1HjIBj0QlGk
xVATEhsIO0iqwwLPkKpL3c6JwV1Z3vcnSP0i+1P8Ebva/3RgTd250YM6DNwN/v5Wsl/aUnVx96RU
lnplA4XEfBLpLncHUEpBdSI5bVPcngSZt0bk3WFo2v5QKVtf7Etqcc/9OqUvtqG0Ef+8sDhh2IJh
jS/1PA+4QgMz4Yg5wJAteml00xVFwgEf70i7f04QhTj/oW7lL+d3ozHwMjuhNj1Qo6UtyZxwamSl
ZJ7kRNUyuZXWeaG7EwACRQL5Pvu2qBRdBE8RXEYt2lYVTfjIjTrHrSZPw7HxY5/bpwjjJ8WmyaOR
Ea0HTt6+Eua3becIxKqx4bgQqnVlekHt/y5+NFSTeZmse/4tDE5gtSrLaYzPaELNeKpN+asblz7C
rAKBwNt3oB931yvO9jH1mzRSaLBmFAWwg555oOB4KJwDcA+20A1pagUHZHIXC67/0OD00y5r/vFh
MsPvQSHfir7omEsTw6Ur0MhPkkmMS73kZ/fR+gqt0hZuIm2so2liAyKrEFmzMCbaBY0i85Ye10DH
k2JqW7rk6zg4vbqnC6Buq37c/MSCGtVF2uhNKAH7qy0libJMJzOykl1rtCkd/JLiIa3oHb4DAanC
P11JlVoqfI3BLqHiiLf+D2qoI3NAAg2D+XD2n41dCKm5TngItTVv1fJMFgsc/veglqbPJl8jJXw9
7EUgKGrXdonwIkD6lQIInJPEH9jwsSje2G8y7g3jMwtQfeblrl57huM/yMWGoMNnvbF8CcMjTZv7
Rb3YyNzizlIrXnc/i9dNFmTnHI/+Tmpz91Y9vLUqDakTc0BkxEio1MY8HMvXCpB/JSEtKOs/+p97
HPrySoTG9PBmQ6druPc43vy4ei78mlpZYmyVCs0lBozcJS7Pvqk0VqYZFV0jFqyUrcijxE30W1UJ
FX7d0G4kS5sROOYNaoeLlKrnE6Z2n8uiGhPFFYBK670napFhUVbhRuVxBwfh29tqGnvEwsAfVzMV
khMxU5TMZsZ9Rb6m9ZKuhjceih117jNxscBzEvlW71J7VIK/0aLJZOoGdFKvv33Gjz7sZV2iyVu4
vjNvWJYUJ0RJsGUyJNfYwvr3ELn1I0c4+YNui4IYcw5DxMbhteGqJsV3QUP3F0JLo8eJdIcPsEeP
sEo7i0dGNp0MlollN8rr/4s79uIgWYgw0zDDBO5Gh5nG9ytEIyWzqvKNoGty13AwJ/XgiVzErsOk
dskmt5V/EpgxgWOmk6yRYKaC/fE0VcUwIZT/ty3F26A8CHgSiQp3JJ5zFTyM4PV5+1A8Q9mMnbg8
czx7jwPoYrMHvX+9sjuLopNRqIM50DD/yKKrbaZctCyJSRTIRPV2jaEDLO653QHN+9MlfN6W4IFL
iXw417hoiu8Z3sAur9x8hH2gxcvPxNGYjYe6tRbE8/qaqUgSBOQZWfyq+g7cq1qUduf51/2AHo/3
hh/3buv/ELlgGjNbiHINHgYu8qLnYp6zCIIyaWJGSb6f6OVig7Syrlt4YTCCxHpHUO8joha1sB7K
VRasC+BwUHidginF36Jk0eMF99Ci6WgsbvYGqK3C2fSPqfbFmXf6tg2PE2Tdfs/geVqbBgO9r7Y3
wQinNSck5YEHXdys1KZFe5d3oanuJWG/rbZKjR+K+jCydUQIIoTmWvTaJiJqz3OsjXZ1aPJAkAVi
mdfHHdDZUDWtYz92/nexgF7EQNOAlXZim57/RmRHxdD8M069MVe6HSAKyNOd7q+GEDO+8aibfIE9
3VK0QBZss0MZYTLMT8GR3pU4swOIacl7ulUMIr0ujv4PMbwbjsuYwn6J/3OjQAeQU1GIupTRFPzp
HthaRj6a2CKWUp5fv5cjAG5mQSDJ8QB+E+2kLEstEn7qaLsU/UswP20eT2WaKTcoxzWXCf4j5ZYm
DA+LjKOcn/J9nbp+IvxZdFxjdByJU8HvXAvhMYQwA7qqbACtPykhuornHacgnjLbp8e9dvIOGrkT
PYjG+ve5UUgEo5fOP59+WpmlQCpZlc2PGXZymbpPEbb4WxlVYyLN7TvrDoqr8Oh0rKdgUeMNMkgi
q8vc5V/dGpJ59VMTsZWPEYdIu55eUcMKN2lVhrKsf2jmhz66MsY0NWtFVYq6kF6fhgD3iiL9yQ5R
zznTcFURbYPwNhPvuCwSgpQ6zmnCFYvN/VfQR7WxF1ZvhqkXKaM5sVY6gF6V0xijT7MPVW2H7daV
yYXHQ3zX/ghulG9FTnMmXFP9eEU0AsdhShVCiQZAk5JLB08ZaGIC0Yx0rCUzwgc+1CNM7R75x/Vy
p/1bTFTgyCkjE8ngsvZ0UZFTwk3XEJy/kKzTZu2p+vJT6YLz7MAsnEpJl7zYC0riO0SYi/2lcAYU
2wzkDHPDH0ABpdjX+n4XWB5XZS+F1axbS0GPpiENttFKeqUgr2AtqxI+zkbJVMnrmfxS4MqJGBlv
LRCDTugVHXMiW5EP00td8K2KCf9oYHGCFcyliwVo9Q25wJuHUhebTwivSEiduNf9Dg3qW189lWVc
TGcrW9KZYBpKK27XaArSEGlYNzD0PIUM1SWcL1xII5rLWOsA6A5Dk/8IoUShGHffDPJQy+WK5d4f
Hs8mJ31dSTU8ntGt6vmlYCWrKCG4PSDpNjI8mQYi8Tmqwo/RDwn2v89w9Eel5SLw7xmsx0eBa+Z8
99EwlaLZz35cXjv4L3qAF5yEYMdfgL7bkiQGmeFcmqcyyDE0v5RhL33kZbH7axtRbbQpVsVgmg3k
u398hXrKKEIiBEmwhpeNCP96Z2Ay258hNdSuiZaQ5ek+0TjN9r/jhbdl+l8UJh1dLB0FLHcHRyiY
2bWnOvvJZgiks9gPy5qaTk+v3ABShorSo5eB9T1rpDXrtKrcBi7tV3hAAhv1Jo0LVh9FIcICRFcK
OI/JkPKaf2tJ/BxSrcldA85pjiilszaXvyNWBMXbm6M2O9XzosnIF2ibj9DuWXC76IKOUVy+V3IS
lfQ1/sRcO4lzWhG9qJdYIAnAzGbdXBvDx0Of+F9IhG2sDbQaNKnDxaRcRPT94KDTK0dyyGiVPqcq
B2H8RCXQa5E/spfQUcanTIMkZsxvvOztfUDiDt73fMpWHklLEN0fKu9tztTtg6tMYT3EQif8MGgR
YpV+XXAtPAIy2N4MG4yVEMYtxPWxeshb0sHRMyMGoCDla94pxFiN0bs6T/NZOvueLOSnb9/Oi/20
yOCUvf2PPZCq7zyFcHgaSemDUruE3jsLtTji0bCNEuMvUETYcJnXpJQutYuojlt8qKyakKUCfZ0Y
hZSZ17ISj3a8C9xk92rjvA++y2dxGJ4BZ+kO1HZsRHS6tq61z5zQoWU9qZG2Fwfe6V3HI1cWYBNu
cvHmiGffyKh3q2i19so3rYEu6LIsVS/UE/GIqMKubB8TErvcMUDUQREMWe7jlM+UznxH3cqJ8gdt
u3mABBxRQquxgUSH3LmaFIajmjCsH9ignrfGulRii1B9V7do6utZB8JmbWEHvNh3vcWm19k/ssnE
ecZrBCJW1fXbO3qsbe2uQ3BKrPV42trtPdNhTS6dseJOJ+att9wIlkffb81DGR/b1BlDbSWjAHPc
brrh8PgHB6hPFVb22TN3LKuBD7RwuROFpTzQOD7EEKxEeBKyNmeemYz0X4U7q5o+c4Ix3ZqMfEuD
cEtXrp1EpwuSvI82f+3WLidqcQMNmJ/qgsBRRB5grsyjbzAvQq1XUoCiYyIFysZNX4cmnPs0RwPG
fv+TUJn2+AXNltmiJmMTdf5YE/K//FkKZ9IFNJ1Gk2QmsH7aQ1++D46bB4rB3n3HH0mVFvbS6qAq
UMlZKzYeURxdy1kFb6joVmHgPI1I7PcthLf691wXMuZ6WxteDVOYQ36ap2pMsbSo58BNWQDgvtGI
YNPKEyUVrXSK4XYbNxTvxMSS9UTODKYvZhMliEwMsLteXvy8lfHikx9Tt341NxZIRHSeDIWgVSod
xlR7QPaRwE9DYl+KaPj2G1Fgn/MgJi+zCmpXAOn3fkJMZ4fzbKQu8jMUjZNBPY76095vICyheyse
RY2X2wx9lXVHYIq53IKiUeSaBjCEn+oQYo2w3xprh6TQBaldRWDhjTsY8Cl94wCq7bl3/5ExsJTK
catPFhn0mCl0lK3niEa5I+g0zqkqGfBu+z02xhAil0STMw8ECLyGPI80Qa20bPZwU2doTUT+izf0
HaS2H0t3dXBl+ohWmsGX1PrUej1PnojeUYlnnd1g+h2+nZUUmZ4cMCPfZqQVXqJU+poF9HEuf5zY
XBym0y62azRUZe3JkqvZcndL6BS7IyPzXEriam1ThXaySuTJwfSI15Tnh0xxpJzeuKhqqpjCPJWp
EuXzyB82209m2YJePeHYq3/QghyzL+Pd1aQno7Gce2rJzhpa+5i2MZIp7VgCeP4kNftRCuwJJjZg
Tfq5POqYNZ2yvEgKU4FdXB9XZamMzGBuSn38T9xppRs9d6oXeNRQtl2f0SRBQ6ErbIKG1Pqa+Jk9
hiLn5oJvQjXfuu2SLx2USP/HF40s61JLnC/k0jbexvJPwj5k7Au5fBE1a4s+j8m6GYr7uVHq826N
eb0mzVmjTS8PN8hd8J9vGOZIRfV7dclHZn2lzIHIpmQX2wk1icvsyiohyL7soS45BGXl9xrWCF6t
Wdyrit7R7X5kKBNofotur/yPXByVIiOU3VmI9z1AdvEypyR41AjEPngU1MJwZar/2IRo1tOWPCZE
Q0icgwaux81SNHiTtEpjafHrNrFU5w8UzU2myEt0RzwzQqW99CGIlzGicw0BZYMcgfWSU/ZouBQ5
0dZIfkCt9Au23fnBLpi/dSc+MqkAdkMW0GWuN3Zv6BbEVZ1lh+awGMgPJR1XBj1tppBwsvsemPnA
XslMHDt1Xl+v9ZkIve1qPjW/IZXEopA2qypRRfgHcWA/3F0r2GVU1Vswh51rte99I8v89nWYDDUJ
I0fa1xVwaY1keyI6cN6MLxOM4lngRsRBkCk7UPYk7D5u6EKfd7re/xTj9DsdG9NPxeMuyU9NcpOM
A058XgoXHK5Cl/RmThtkMTcAjsmlmhM2LDlUKBb8oFy/GiIXl/9bWu/K6rde1LMpEoEYSCOMKkLN
2eXQ9SHwNGO+jWQt69Lrc/QrM37YA1UWA2AlGD5zod7rwd52m82bndaZFCkZ0ii+sD9J4YS5EDQt
S+htQje46O6hj2jncMDepFnAIVroyELgsC+VI0KYrGaYbmcbRuGUfsUknlZZS6Qs5ysJBWDaTKHf
lu72dJetf30hIda17iEjeuvWGaruSOIGUT3zpB1Dn13bKG72NcZFXP6qY2BbQTOPSBMkPMXWnulF
LudRoxLae0MpTyfB5TaJ7WdezxI9BgV9IBN4+iQsF6QkDSOl2hj0wugNIdcDyu6/gbtDKQAniISe
9n3owrKjfViOx/Tp70p7tTWOOoTEeQ9yCsXSaN4o8RRoH/PE+mCkKoYkqXlEvEfQ1fq89QBRGDKc
3txBOF2ElokUdhb5v+Y6ezfrKIeBdY472hbf86WiMyeD41TP2hroz5NkCWyBtvsdtfeuEyn10JqR
NUvTDcILLaJOkM/WX09LUps1y1RwYEioyeL3NETOgXc9rNmz3jB3MOoyqsf2kU92e8ml7ZWeyiHh
GGXCa6k+SJb8ZUrUIfTQmvuRL0d+5+k1LE4RfGV1ORooqW3SOVTyJoa5evZEPsw037SgP6R3N4kN
tBhmUYh0uP17pDXqFWm5O2dLC+vNFQrB22k3EYPeQukiHxvs2ZfbESw/8Oy0WaJkPRh00YpdEjqr
iSUKw2sWbgoqbKSY9w4ZQVfI0/V6W3VYACEfmI5dSnGIzver0ytMhDrsISbOVE7Ei6kQE6Nsztzi
vuBm8ZYR/IWNtqVN//dYM3JOaOBYH0jYVfHgQFqHxsL1XYiBcGCLir0+OOIGJ07vUrhVgN6jMB0G
2mzK2Y3o33WtrBMTSTW/0Odeev2Q+LQ+YF0uDo4GY4MbHLGJ16gqwiaYzYOCanLkoazrL5SODKhT
Zbiulm99hmI8UXqdBrdHAUjd/xknn7XHZf31DdwseEe6gwNA7O57bhIpa33Zx9czE7iV6+7lnn3k
mu4k0qtNgqvUZ/+tEJhHhyhjcSsgDPCeX9c7PkegYyOPN+haVOtVj3a0Yn4u0cILwfm/l63F2KHL
KIX3kUmUherAbgPOCOY4us3KUyXwO9y68SZFgKmipmtN+flPGRB3aV3h3uU6h2CCGJIsma3KkPPH
R47pNbxjkT7p5saRQ0GZoGhS451s27aiGkjtjLWupg2o/9+O5AUwR7fbWwb5RM07g4ziHMea/SOC
9j+GJZbrZco44RWZ7ZgtmFA/d4iEQQ3sZph5qShV98mE+99fTK2YyX+3Xd1FKdzJyxnpo5b5xlK6
Si2o8HxaY0DStWEX9xipmQrhQ5EOhg3PwA/wZZmxVEb4aRKFLp+a3yd1AvSOvg0sfOiLxs4qIBA1
/CWkB8nS1Wvr0ERB36uqtGUt+QY8DAnzYpAaqV5T1fAeoaufx83DrSBxWxkovZtAU25SCqbMvj/6
TZBIrpKxcu3M66R7Bqt3Aildo4JyEdL2hEudfnn9h+tPDizDxDSXqYmSXrQ36eTJTMp5/ub+a8PN
mkHtniKwo0ojbJcTUwMGdLFaS0X6GdR/tLPl03CI/uBUtfIYGy7NM2nt/DOQyuaiGWv35QZ592Jf
7eiHabtAxhS3q5u/AYxjOfdcJHpe+avEH5mr+3UoXUCtQuKSzHJ2c7PAvosebsj/Z9LosbH0vgWO
srmrFqUcx9yOAaZ+YHgEyD0Mpq0ZQ3Ou2WoDSZRWldBUHoMpIeHTTwEeQlxIk8ymUfLmg+/tePD7
q/95zCI6AsG+XjzCjTREoJ2DLRV3AhVlzRhJoQSWwCsvu98siZ1ofJpca9hiBJDRQpogNr9k2Y2v
l1gP+nUwkFGLwXSBTJ67SGaQ+acVT+N2NZ8nhifiogl98LFal71HxmMz+C8vzWBF8lCjS2HZ/W7u
0naGPbIFM15H34AMIojeuMQhr5YgNRljoFBD0T6jxJFDzEg/R4wfSJ6ZFrxIPmbjqqW7ATrtVM9m
1E6+UAFvb/cbRWtW7RWW2oPT83WeVqrukzJVY1MV5p8HNQz3JGRUMR0teQW91R6KYRTbysT/39MY
3w+q/NnB38aRfVX+Z14eMhqObHQDbLbSxt3vfTIvZv4sCG/XyTxI+5finfGcfvTzM/94BpagbFal
kF2yrnZVcSX6WcPcYE7sKHC1oMaabshyNyPMggWC0vV3oPUbSxUVk5aeb4xjk09sXYGT2NR/Sg+g
hQk5iEQW1kenFib/3phyZ3ufIu9bcppTyHhIKw4qwfWmSQmF44nVDJrKXod1ZNKx91LnJmpmrtht
voMdveTUpuoRUm8T6FzFyL+5gbTycj0EX78wiRoZeXVw+LI0pnQ3CJsB+DaTVDTNyQQ5dQApEYu3
++t4RiWyeFRNp/bBSBV3aJB4YB0TX63rpymfIGH/EKfou+fjGE/go8KDpf3WlCsto++QmF43ZALR
MI9MitaxJuPf7Da0oEgxODzfV1I1HZraCNX35Yixo9f5wramcc6i/vCp2akyoU3YP4ZL87AWOeP2
EdMns4HJNxprGp1WwG/PskpgOJhwkT3wKkNFUbEfBTsRIrkYKvYNrZOhRRkMmHlhidZ+YXoDJ0kF
Gwmd3VqfbZGRUmRe13PHJceKtKEwRZE+rwlujPB72bap+GJYWOmTO06zEY9OCIoo/bx56DNEJKhj
nTsHPsumih8G9iYx0QljM1p5AHa6ywidGowyrQynoe8hq4VFbcngBHAFI3tb7eB2qCZwfsg51yrl
3evNzDKhVi/oCSxtH1XKcMvE42Vf3ixABYr1eEm1phAzWL0S9QXCkLtrpvqIA04oa1bm6h2+OD6G
CuIbhCkg7ouo6Gsop8d0qO+skS4R51OGaWGfzpssM5tbvAgyOR5NqbWbeVsSnO7Y5lQGNCOCv4IL
EXxI7WZOWJU+9mq39OjVJ7eHDJPIqqzWRq/If5/u0x5vfDUXjtiRrLhz3RsAuqXW3h4UblXrsQeM
adL8NsTmmciNJzzp5bS8HS/mcijEmoU6YGLCbbYimftr6YJYjLoOQy0El1dMLU1uMlfD55cn8Adp
f7gtGJ25nOr2+bTuKAmEvVfHzDrCfjU+P8ci0KsSJdRukhClI3keSE6at0kalq3SGjdYUSWyj+fH
AbnoMC7MthOtySxaUUCje3Jj3w+aIpLZo7r/tWoI3UJ6sTbt8f3e9vvLIdq0c6Yjv395kbWxW48q
fTXKvRVOCVSukBpn7heA50a/0B2QFhaV9/UZdtFzpb6Z0ZkKUhnpLkbouRRUjLDyBYCp1uWInb14
yJStii6KzbFC09DB84Ds1+zCWDYu+rcty5+tj8gUjsAi8a9xxOUQoV9K1CDLMukVD1bR1QM/pjbH
G6qLPCRRVHKm0WIre1GTNYi9ppDR60PkKK45+l5XIQf1Ei3XnJ9z+DodPcLyvZa/mTDE8FkqdiHg
pm8BSvQuNNe6ubrp9+goeHf6bRXSFXeK8ijObtlSr/F3T9mTISfdLsGjvEGi+liTUj3E5D3dIU7x
22Ra4sVHy/9PUNAIsKq0YOWMBbVvPnf0u/F+SqGVJ9UoB0Fv3Xb3asYv2R0URDWJwdHGuywG5n8h
o56zkQ47fSdngChOopTMxz0+Wn9s5m7a3nAJU2Hq2BV3ROb0uxmKRXmuXZUUVSmoLtHvu0dpBVlL
QapN7W16aAc3RkKKE67mJIzTirfICc+zuK7jcU3G0ds9B4Jnlj0BYReSAaGAphAdF+boDOLnTweg
TpHQ70Vwb5Vui10piom9Hp+CFN9ct/ru6WUAElOxmsvp1zwM3yaDjOjmEr3B49zRQFDI78V/ww97
lrfiTjQAdR8k+t0JKAXsCxsTKEChgAYPNZqpXER2EjXS2LNz06icenNxwLL1YH11TpQkwnkhuYMn
7/lI/z5x9ZJQFgF92n1ycITqDSFx6lDFAVVbZY5O+8HIsDxb+aJYfHSX5/KCWh+ch1sRUAfodf40
vtGcBwLZsZNyS9CCKdZOZOO+HrI9iZgcAAldC3VkJtxZZFjJ9dcX775jpF1jG5LEmH5TXhzF05Ra
/Iv8QoLtmJEpSCIoFFp9oFoIIV9hE58DoFbLOWTEjk7pz4W2L80QnR8mguArzNulP3cfBSAOu0q0
LVK6eAyfKIVph5zsnA+a2pU4qq9LZMi51Kw4tDa/uzBYpBxwpuNG0erBIWUCjZYrDsTbR1OKN2Kc
4kL0lqKEPbzpreSr6BvEzkOwUoicLs30tmjifJj6cpxLYOntYpYnjtqWn/Ix6k8IbcQbl10rk7XH
iNgQPjiD/ooXfhlEayGxJUBwzcsKpmRXMXbmb5blSDL7mPdnBIPaIsIS4OyUkj9+AafWynZjeobb
F4JT6CI091ubjsmh5VH5IIfIu3kKKVP4e3ON0J3hWLJVx+HIbfjf18yZp8r5E08nZyemCupAfaLW
nixD77rrrX0xnD8tMwTkAm55B0N4HzknFVU7c+SOg0dVA7mArpxtgkcAD3fJfgTze3WRBMmQBd1R
HXE7JTs79PA3b8hOeQeZ26vRkf88M1GlwrR7XWp+N/YrIfEs7ZruNwooP8mB4iPoVtFh/EYsF+N9
ATdJ6NfedbfB7aFE+7oFXqd3gBdY3uxWnvoZCku35kwoHJSa2m4QFg8t90FYUlB9m8RTpiKBRG73
6v2a6QmMwEGQDvtS7wSgYwbPmihtYkLXvCHyxnkPGj6A1m8rT2z5wyF/Y+xhfOpyLrOG9pE0Hz2U
DvFwIlH4n9KczfMSfA9YsY6sc5qhqWQEUFiUnvH2abT5nlDJX0lctGcxGXV3hL7wnn6dH7nVpebt
nIhDOZSax+CVHGkunoDhZYiScbkVm8c6twmkKmnnDt0fwb0vxAWbLQV3wJLzqajR+25++RkJ15xC
ImPzbvAefWtmgu7c0uLDENwyvMA5/vPrKkUeWO7XQLz8tvI+qdU9m9vJfUgrZqk45KWtg5FowLLp
nSQ7WtHqQbVb7t1Al5jQpNG8NX58So7kYB/a7YP4GVCm9in28VHLYQWMIjPeVJGzUNklUMbefdyT
SFH2E6uBPATZxqm8lOTYlDyNpzGz1UppKUfTvP+Yh4DFox7gdDY9kTXt4kZKMFrw8AuaxoXPlSrL
i5bHOFUdHwoi08kyDHX2gZYyo4ucBA2vEqXL9w0wvl25mKKBnMMUmXUUP+t0Wo9+dMyOk+I7QQIc
3ITm86GnbuyUG4RFImkPYHM9h55v7wKdp9Cb6WhsJW4LMe1e6sfOrZgBvSEgCDBravGvw1dIVpq+
gvsRJAwlKJQ5Rm+EZa8awfp+/34OWBcUz04dd+BO55rtOMKRSdA09TMVdAN0+JBdmqX3o19EtFz9
87juQxXdloom+Wg73+bf73RFb8s1Fc7tGZqK5gHQhS4a6NZZeAGTlr2BasE4/gSpUTI3Es9Y66qK
QiqLsMZacpqlaHzhb91JgA7pIG+U4nh57s2ZAlKYgRYPAXaIzEoBsJ6sUn0DdvCLEotB/rivSiSL
4Y3ABI7qQ73Ne4bkTMME5zfeVNfXIV2USxR0Lu4eT8JNKSlTMsWYgOHwt41Y15Pr+wP/Smb1RNSS
O+kQsPDwzPbzI+FZv7Cc7Lzewe1WliHKiCLbGeBPSGFDidIR8DSqjw2CqqybtjrWdcTOS9unpjP3
1h+R0r8e1boQ5uHEXmYKs8Ot4k6NUGE8Usteca7uTtkYY3dQCdc9ECflG+ZZRrLchsLWVRVluufj
OJvVa16oAme42wNXUDmi8hQQgFmD5kwqJBsNtIDSeXVVp6225DMtYiec7yk91DpDQzfgpShrzI2p
Gc4R4vAI1BC3bkhYuF47g2AOFn4KQ7mE5x48wA3AJv4VyGykNQb2RbmO12l8FdpkFblBIXwBfPj2
cjd6R1y7Q/VlghqnY2WhZze/4qeLUCrhILdkOkngxMvAZ9COzGP0GrwqOIjutZUq48nrCn9h2rLc
iem5rWef4eWYB48na9AEoxj0kxrX6dztTFs4lkKk2YHgila0wbiFY3ISpMs5sOQ40lao9wxWnuoM
f2oos1rHUSUEAQAF2jHn+XyxKARXOnfHoWNzvYOhqmHhJCaPcMZ8c+BppLWAkTucRQLzijjW9boF
JY2GPeeW1d63bCLdQfJ1N9W4RSOVOf+7pTtlQnuAQtR1YNkVGiBTzD54dc6ASoiPiRwzbSE4jjRX
kkWsI2al4xg/UPb76gZBumIfOXR7gJ6920xZOBLVQM43PWw7NYBWCQv630UBNdv/aVz9hojEncga
dC68RJQyrjIXHeSyb+MDIG1tTKdlZV4R68SZtEoMWRLrTx+hjUBquej2GDqidM9l37QOGBrQnJP0
hIaYQJij/inJAEjs6SA1S73JyNKM5jmsGZqjaVFtLj+XgR3zND9De+OUTwpoJF+FvsJvUUXcnHL2
h6WLgXCy1eK34oE4iYt0AUKAD9PZdXsNm/FRspiLaDbdHL+Ggv5ILBuS4nMjrlaGgOmonRgmaVWc
CWIHU9ytBDUp64m4XOeZsLW4pOQmnYbvAib05JY5YxIhlzuY0oU+4jIV+cweRxSjWwGTcHdb7mth
ICNr4tMbj3XycyghXwe7UYDuCG7PRpyCx2EaToCIK0LagZ0qCcFY/9wwEZXZbS0WbXCVb9YnQ2AW
MayzI3gRXSkIHn+6bCThfe5H86oyX1ReqA4vAHk/uFtAJQgOXCK8wbP+U94wOBFPOkMaiBVnqo16
/FHCFnRHrGz5e1D3BqrIEyYdJ2PeWKQba5eTTVL9UuPqI++8RdpR/DQ42dbNWhq9OSn94/zTaQEn
W54+QalbP1K2fN7rxuULDHUfOJDLJkZZUFlEQuojf4OWsfuemL0VOqjyZZTJoaf2/fLgrRFD+MVl
X9OZZbkDwBc9bX/E84YqvUF280WOv0slcbsDLaJKxtz2j6U4dRgFLorTyBINMLNJ8pTYJ/2u2LCw
TooQRAnd/mg4akSuKoqE1XhAQed2jh6tS6dncCCLKC9WdIULPRajRTAMnS2oR0kH+ob5VNbqIXGu
J1C63dGISEVcqGlKmpWRMaqW2pI7/2EoqQ4FoPZS9LbHaJTklPooU/wi9p6fiLo4nfoIzHIXJn2Y
G7Hyg6mGe7ZFChwcCFH/Kn1eYaC4BrBgn4ThOfGpr/t+BU8mYxdfcij++Stwj72be3ZYqZC2DfVl
H1c/pi696aOTTxibMr95d7Zyl6dl33L3/w5z01OEp0oGRd9boQKdaQNViBg4ZdsyKEtZH7TXsDwm
Qah4fwJD1ZuL8JSYOFyd+I841SZpXCE4UJxsyNlsuatOgy+aSlhTa7z0DT7OwirFjakJcIa9WtJP
9R5uFcjc8WRUZvnJ8Txd1v/+vNNzSuOkezO9LwPwRWt0xfELaIQ0KXvIqyGIrWx09YYJ/r6+mXkw
5eSfljKnGcdeBHvjluWHrMR6H0b7G2xyfPclgOZaMwTtJTGXJMV1pVlusvCNKtQeX83dhVAXLu2r
Y2W3tMjaDcYO9hFE7XWfDLZkzEsgXoHqtfViju6+nwYn4vf1SB+2RYIwE4bMeg33jo9TEOmE60e1
uqswceKu8MGHrdfc2AV2I9FGUgrmx7iBtBT/OAJKk/yty/4acIDj7PnDzxH5ffidrIe8zTdesFpC
Lub8Vl8UNPm/DgSwjdcWV1UjBf5AuGmtqzsKmuyjzJy+Cp+FwuU4iz0q0UsG7bAdENffsShyNDuh
qL8lhuAteJATsJBfj5tgobZT+CAQaoD60zrzqhZfZSneEpBKpce5FYfSJIHuIwXX+h2UEhBjMEki
hoVdkhnGjDIRLbtW7i4ILb+HqOAaxEQo4HGcYY9fhO3tO5r9v45f459QaO1fbBUg7A9faUtHkFjt
LxXJ0bWKBDfnpWL7rugFebv6JFoFPPtRjU9yOWYWHHD2MPkfXFHAE6mZu2678btsTpdBh6l31zU3
srH1vUv4EaQYhmLZbKQK7uqWE2KyuVTeQxAzIoWcCEIR2UJQ6dc5sOgGN/8m+CldZ/m9Q1cgHJ6O
G5mAwU53FJlxGDf9iAYp6uMRJ7Xc89V+/5GEK1cf4wdSOHINymAgHkjsYlHbLdW1BUxraW462t3G
PGQdKZyCldPc+kKtO4YwTPiPtPagWdPTXaoC4iIozGXbqhBaraNRksr3jeojiw5VH/4itUgrPEvj
0h2G0/WSKjkWCCcVm0ZSQ+0zgGDbslp9dbsPJdYFJf6vpKvNqyT6uDhIFWdUADBTJ/Qo6fQ8BGbQ
/aX/hU/soH7hFjVJPNq3XpsiEo4aJVEDpcLLvvSueHChxwH9bRU1+gqCfVZesMPDPuSw4gE84InP
H4w38/DLyMNMFqixoL58RFu69UkrD4PZrQsiv9ta19slPwzXfQUYgflYMz183Qesz4BfPXMtMnc2
wmJYB/CfZYzoBKJilec1FBldy8QmY73PI4KCzfe3lX3yuzGzS87Zki1TcTdWP1GpMj1tuWkJ2hG8
KNOBSDi0IPhESbC86sAps60hgQvDwOwQQ7nx8WalCi6ehYXe7v6/AUek65spWdomHfnDb5UDVqVg
6Fim39xotH0bcKQy1TYSOnZ6bFgjqTbuLYh8MUByxhnVkr4/RGsgXfV/0pO/AyKi2d8D62IDJX+o
3Rhz5BmbT2zHIYWKZDiJ1WOuz6ehqWK+e6oukUtV/7G7vzHnpgnIVsJkNhQloCx5rPNKOVnQPjbb
2l5HYu9fInuaV0PV2nB66bDj4tJ044F7gxbgLcs5zPVcgD6AVNcu+PjurXmzraNimaAHTn1iLMdh
+L2WVA5ErrX7lmPIJotw/XMYazkKmn4tr+UdDiqfqrVlOjIAHtQgF4yRqXNkPI3/aG4sTls/8n4f
PubPpbQrG/oBJ3KHyhSA0Y2tKHMI5roZxyeVF9gVKzz5/tav7tZW1neRK36N6YH54dEOucHJ+n66
41kTNf2OHCCN/gnK60ogku+mEa9d8JkVnjRTJJZiFi4dSOGNgkbhAW63AUMtsjkGWf+uK2J7jaxO
7AyZK7IJvkz0yqbRBvjZpCsCIgMXvcjBVFWrP9RDpZLVzPPz2FY0RcjpRtBdva1oBu/OMFaRadDy
ilTQRsdRXQ1bj1VbDt5USgul487kNF4zYXE6IC369D6tbMUe8BSLiZ+9t3d9k2ZBU2d2obnVM0b+
opVmGlFeHCB6kSrrCk+zvlOcOGk3+vuQm3S1kSEw1CMhsTOWR6kyeft7sME54I+0hmb6eUBqLxh2
QAqQciLyK9wmUMjDfyjTbNxJWeASxwrMEVLvOfwvVZENqiizx0sbloV7rLC4W4A46OA67la39a4H
9xXls1XaoDWwIFywdZkfk+w41QtLMghNi9NOlqwn56ZAxWJltQLfn2sAN1oPnA35uJkQRbGz+SLc
xvFuRWnPN5zKtxa3B6phEBZrg3+vXDoTCpi3rn3TEa8HEawQJ2wJfkI2kBCbVP22k8VHweaShTSP
cMUTJY/Qes1JRYhtbkpNDW8pzbY+g3FC5WtHsgATNKzSE/sJ6cXWbLCf0u5i+pXVoF/3KHtBkBXx
9+d7IDFGaLP8Fhc3mhCSfOHJhgNj/E3+YhUo/7X5So86dgzWr4XovC9Cq9J89hPGsmZpcKXO3d4l
zx5yWLohGa1AtSqCwiXwUegRqQFDouiL/RkG1fZZ/ZJzOrIaQ1m83Qq7DiA1kHhlD82sinSTQvtV
ec2oaOkGcSzEjOqNE/BwGDa/gsBV1FxOGrTPG3gW7euLxGQ5xASNWT/f8mBaEd1crrD9V54Kfg78
n/ygwwZ/Yp5+nOh8yr13aMw6r5ZsZvlatIqBp7/yNbKlsjhhVjsRTY+C4wL7Ha6r8uLnNaC21iub
DOQeqES50ynRqTMUh0+mTTTIBKlqYVXDnvBYiTJu67v25PqDrawV9DjT8mzxv8l50kp/Unch/EW7
Nf5+0e2pVseKBlIY2xqVXH44ErOhX4LWFfmJ7SksaJQBq7HsFXAS9on2IiL3jE9Yi0G6o2bqhcwT
PRbKi6r2q4YBnrapkghnwvrOuFZo9u7X1lM2pZSE5UCFHY1UmoYQ2PjXv09mPkT+2akE2BHTcP9Q
qTqrc2+FY3pH3ZmK60QFrvjT/g/Ry71b/cfSG7bCBilOb5MRjDsCBKnJ8cjP25elaqSH5UJVi9Oa
zEh/+C2i/wDwOsIR7u5UziuXcpQqf/18LsgFuTvgpH0LCJga5zX2RjXliONOGDFwqIbYBxCCRjuY
bhLdRR1oVfUGzWzgyqQsx7Bn5ludpZMU4PEEbejLN1hl+pOynrUCSKQ7oVOPP5em0Z2tOZbNs+15
fdFkTbwLIHZGQ11Rqisrsw8h9XD3VDwuET5dlUME15vcqIo+pheQN8xHPunhn13PsbPx1TznItpO
Qxk24CymE1s11tsLEiEBdymS7LhyUov/sYQJyQ4F6L662s55rCHDeFRpMVK2tsYNJ6HktT8dtIX/
YQ6ve4ycY8H06epESmtP5+4w/WcdFwjVkR+qTYd8XJpwtJy1ZmYQf7vgthrKSivPZkGBGycR3WVD
a1w6nId6RaaITpo5QNWsPjBk7wRJqSQtYk+zceNUGwuPgxVAIOeqNhJnGucRiOx0qUqQywsmKmt+
wwq9ZYwv20ztBNoUeMLqGPEx5z8QKMXChISX1fmDf/oEJQswyr4wmUEA86ci7JFgqW45m5qy/0Jk
thBalCNx2Q0iiV3JcvvG3LYE+w/5+zm3js7qIqGinLXGPhoL7vARXi4aJOBoePdmP7LN6asphkBN
KFLfM7TsKZsWLWHglrUtwNaDDDsVkYJZoaM8dzG+13+8Bhmu0ObBqKf44rIQ6x54Pwaf4BHmSvQF
CMf2CUYdUSHxZN9gxS2icQTGMauTRkSHJFr+xKDyOeT3cAO+ZpHS4sIrD67KW1+fzq0CddjxD7VL
WQqiuvdA9S1E9q7XIY1ThNHWgxoDUa+Vt/ETwYWTtEE71neuFJcqtLgtJxb/mutL2WGhYvhagApJ
MwbCsnmNqfFsxSPyWXi8KHyteYjRiZOAl5rMu65aQL5JIR4l2zNWSJp88jF+De/ylgmbtXMJj5Qr
JvtSNGOuf6M2z4xCMGysHqqPyMR7jAf3y0/H6XShYQacqh3rNyGKQ8AKLEVmUP0A78Ohw6elQFUN
TsHX9XbgClhBZpiy6B827i/iTF9IQvetygIei3kVolw/8vsBzyWNtL0/yU7SySPVt7nB5r6UZCZC
7WRkPFAPP5Y1djrLqLHSuB8lwu6JhvNDOdFdj2UOY5dhLyjyuqszRjFYr1YT162Lt/GluHVAyhN2
ZJnBmoD0INZl+bh/YkOwuriL7KiBtERBwPyGveuEhcM6CeSf97QhRfMxC0DJmK1uku/fyor9JYqf
qFi5BcvoLuZZ8vqYegGJ3zS1/3dMyoKVEfuSt/HNfKRjDWjetkh92AWdu/7LkhZlsatoHQ5sEvIp
DDHTXlza8scdPQxchKXLVftHnB2KrCMJf+fwnnTByN2N/ZdF15hbWv3y9H5i0UnBU5r5dCt0XD3M
zn17VhJIoD1Nt8k+YBG2OwpCMqphB1BfhJA9dQ6KspNkoorjfkJmSuBb608XITVItS0O7qKtKn8x
JvWiXiYHnvfmLsBB2IP7dAtR5eHnDxYQI+buzWxY0hAwA43ZMZmsVKJMwydl67N2RWpI6L0gCKu1
j2J09fpIQZWs+A/msJSDctv9V101lmJyHRz/D90W69HFAUq/rkqMJPZ4EQG98+jd+4fu7BSE2ACo
3LLS49ZNQIDyC9jTlYkl+5czAieQbk9Z12HtS/NNTpQDKApNsfXoa+lGS9paoUsyg/jaOQDtmOhb
mpgPu7YwYHEqILW+8oW42R7j9ttcyF1LgzjIDL2+A7Z+3sN6D6ybiRebo8Vkyka2kTEk2H80W15B
bS2nk+nxvAFp6x6Am/aqArsvSGDSkZ7+xMYEHGDZlXsFMfB7qInExXow0g/LjX0TjWiGQPTmYZv8
cenAWyOzSAqeScuJCiRKSJFPmCDaMx3mTCjK6LT//uVfXumPV9W3ZDEHahV2PPX4VNwcwHpovZxF
QPSai5McaqzaEdR3mPn8ATOV2srpFMkHRefZKI465MW7WHpTHz9V7xJtVkJXBy117VLPN8t7OETX
fPvLZcj51Nz9qiXW5fCGOnZxre7a2Etm3fkTjTW7cHTnG6t4jodBRPVY8HsuIM+G0T9k/3PS6JfR
vu8CZsElrybM26MJ5hXc24tBY4IkgNGpeeaTYuizj4Qsl9vd8SNucA7EqhLCK7FvmsGv4MTo8DGq
fLJUvpciGlZi1tJ3+z7tYVemahkHzWHpjtA0BryAhQURbkqNVzfbCD1WtDi/I973TgJ3+5rsxlPJ
zxUjKQ5m/hOcXTMUREBBLb/AeKfjJigJcHxfq9KQNJfzaguJmsIuQ2iVxRAWi9xyOgL63uJbXL0I
7zvuEqpOGv4wuMgKa/YGOnpTlcHV+wZJcCcpK9m55XLSmGOv1tiuuBDX1k3i27m0qBOaqQvAn4kz
1XJDEAMAm10Lcm+V6csQTxItmWJhSqLYTT3G+hPcJPogLhgtQK2ayoKSjkksK31wV29pio/KBYXT
/2EHVBTwohhEyzMs19urh48MQVYdzVbQNTkKxckupKh9fyPEHagsJCv5U7ppbS/XuL9A3ny46sXY
kiVrb98c3kJiOvFq/Xq2cOswbNC1J8C6oAb2WWCk1XaBbUJhHb9ncouGpcRuOMqJkN1VaKq3MjKN
tjtTP5g+nWY0FJxDv22wpj1/BuLy5JqbeVIcchl+9EcKAKIGfuvlWEELMbWXiiXeo0WvF6zDdjTt
io+jCGOPPWoUSWZWih1v2Oq51+YZFi08rrhIIHFPs4LVUyaG/WrSlcZLl45Ve8aGWIM7DYM5SYR7
Y/tAlBYIoTuNKRSFcs5QBUzc4fsa9kv5UGeMCZnZJi/NuDRbZes+JB4gRXfoYORvip0XIN/jK3iw
7KJid9YaIL7+c9xcFY4kvyt3F7wOFkpW3RGlCEz0jVwy6VLOmFhvUL+ZecuebyxI5srH1l4w4c5G
8neDE15IWCuh3RnFPbjSrSDAs5aLgSfVSkTy0tPaqz7S1ONTWbXmc23fAJfmsZl8m3z0bG4vscr0
6Sb8r/oik/wOupOOUkPGzi3v2Y7r3uMeiWkhpIDAPYjIUB/HLrxkrXyp8c1o1eWacsOjIGGsaxhH
tmeQhCLSqXa4AXYW6SKfizzESvQc/vO7z/xMC44sGqncNTlZAfmXpFYJCY3mrn8/kSV6sMz/TXaQ
vQMbYQpTIRCAy7U/fcwepzjZZCYyuCdSHGsOL0fLDLfB74byhoPINeAnfsU+a4NDKXZ/2trjQbFa
waGg5u726Y2cJuRC9ftUV/PZFSbnu5bNcZOuxDzFDNoO98NhOoao8GZve2JMVYv3ppyfM6HLXdz/
SHrmN5LMKEam370JfzpAq1iJmyUt2rmZWIP2/V1lS4wsFQ03t5wH86UpskfJAF6StaZWqAqALst5
mZNoRokl0ukcCRUMMB73buf+A06rlfwiSX7PLNbMnAK+RuZb0Y1SnumXgg8sE4Kv/H1PoUB6qoVZ
cSiCMZNio8HBYRZPTP2ChFGLQvH7EQBxERX5FP8IWBYWNEp2azyRbUXOroWybNO3htkhmOKKwLXl
ElLp8UCqudFpalGFx2uFUce0QHYgKVf2/eUeeBIoFsBDX0DJG2LrsDZHr9cvXunwIybeGQuVhKoT
QOrnfhERb/rsJ2qAkN/GE8N5tGHlSRes12Y2GhXwHWu5Ut5Wacwz+jXv0mhUS95c7TRYUUCp8oUP
7I3qpAbn7yQ/2iil9sub3yHFxdDDa183O5qZWpWcmj1EKqz79ImS5VLs0nO25A1jI0J1rFO1zrSH
PBmjzRO8jJL1r3fey11QzIbnX7u27jfg3Cx6Z+YkLOllbqBeIn9xDM9Fu22a7SPeSV1oSXVt9gHU
vmp0NqOZ4r366HGRb0e+eLLcxMrBy06DN6EFiDemLvrrs34G/klpxNR9BsFEFjXKwRes+S1/4+kR
Vu+OPOgQPgraXmysIa+NYZR5QNanvXIxQJcEX+oofAPAt7vG/UwCBSAci3gLGKHPti/VKbattsvM
zdQ+pDbryCPoV+4LBMCpptLGfueOkvwrIlA7KQejIO8QlMyU5S2xes4P8MyXYQjBsCsjoUMIdiK4
vkDOuba6sPAP9wqypwMhTjZvnccSrhGDgosRNFgPikUEmI7vbtVdNVFTV4XBH5JyglMOkY0GVTXy
YBLNak/vyOcNWQdbCwUxW8gJ4lh//BdBWVNxiLDf80X/Kw/ayXRbTl4mswjXg46Oj2g2vCkfGj0H
jA/7Rf/2ymhU/jYKHv0PIsm2vmnRiOXXPEDRlAiUe+Lp3lcHYpZcWJaTkXs4MfW9atev3xSpgWrJ
6oD7g9t1LCcQXsXHDFijJsXMzJpMzHv+tsvoQBmTrO1p2re/aVn36SRtc1mXsWiBd6HY5V4wm2vu
MPqVfmGuRB2aHbUqRmZ+sH5cLT5FioZS+zw3ZL+kF1C+tged2JhxyHkKNrnJcGZDJxfz7B77aI9s
G3CwaRAcJvXqOd4yxgVyB2TWEedlr0O8NU84Euz6FiRqnClnxZ+5fj9o1ktj9ZqfaV/bN9AFcscK
rfUGy3CffKwUjJe4tek1r56YNIZTpXhjLdgFlS3VnBzTwbItNsk4gU/BSE7k20o3t53/bsFflzSe
lBnamR5l/UBFOxmZ+XU3+xWPu8uahBBqTyrTdx2utX9ztAIgeE1FTWpCsZs8Ezmfvgk/uW2ui6on
jU9bk5P2WBMuRkRckvJWN59l0gH6MdszmOxj8Y4xKYSgRB/vSwKhd22QIeSKHfdd+DdGhnuROynU
7IUL5jKtPe+AYzwNekeEBnRciB7W1AFGWPw5WJP1PPP80Si16HrnEqlOPeDlHg3joo93V1cfLpli
VUfWXnOObE8tKS/qr1l73JYSUNoa574iCyhpWRSaxT2SRDhRrzlEteGuSugvUsgGDJYKNNzBFi07
fZhedsf3SBRiLu+ZaPXkTDSGkfuONdq58wdSdW7KpyjxhRdS/N0cutEO2qp83+9y12ZEGwfSzbYh
kTbjbGxafCvN28H9/hB3lhSSTLSs3DM1SE68KVdERDKx7tJAH3WhIRiXQo7NHspIp3qedEjp8fn4
Vb5NHm6U8RBjweMGVCEdpmTusDW+SN2YGeLNoTSeVSfM7GDxOZcmR3UtAStM9ArQ+npI83q40REQ
w+9mhTwV72jvpzfqD1LSUx070FNeJNNrcK6bzLWR6r9pEKqnh3wQXpEF+76J5qlxXk+gEeAkvkyl
xyOGnu5pd2sUGX8FIyAG32MhmiiuVfhatBo4MhQ1Fnr92fT+mjaBgB88sIYpFZECZLuPiLndkZ+v
PZH6aNP9e4YK7hqrdXNslvL83YZJQYjTKhYoprjVvVBKXoJIhVZgmS3Ol8wwtknZeEdjEWHal5t9
bepgXee7LCo1RyOBl9k/bSojxwg+yi3a6yG8Jrn0vmEHv3iWj1lqMy2UV72HKN3qgyR51J01DoGK
bO78dV0jE6TXGElJY/4yWA2nhEW+IR2FCR9Mm8wTKUPlHyp5c6BmTsdxTsUBtAEpqkwSD8wXEFD2
iUoc9VjnNbQD90QdLcnQsYGVuvYrcfTaRYqwL+SWDPVJXLzjc6fZsQ09eWx7fqul7rmmL7oBuzF7
6zpIbRnbwklZFbSJHGiVyv/FEQBIzXB9oegtdIwAVvr+FUDi6wb8JjRGzlw1Yd3/jM00YLcFVTYL
q3xFrx8jgAhbRXzSK4UQe+3+9ni9Ydzu9iBuinKpKKqQqx3dyC9RmEvIfrgxpzhreMR14lyAjqyQ
TSveeiD6xYBj8o2q9k7v6FuDolC9LJM+vCykhetmk2mw0/QeP/BKmzXrOWzJP75SzLVWnfHU3unA
EIPRyNm1vlZFNjy2mSNLFGnJ/4bduEYvLGlT6OP6VnLy8ZP8E/irrUfrRRdm+y9SfhtZ/UvTOJbG
kGZ2n6Kgzr/Urls0S19vt0AzXbti29TfQrAdK1Kb7FTeGsN6zMc6EhjHsWNdMuSXp1Mj5wfMZQQn
tKs+kqep+hJgXGq+zp5l/BIEzzfhv0p44DL4ycWZSobcRKxibdM9IoHhsmBKucsakG91qr9JkLBB
vSM7y4H6L/cG/UF0zCXgUdB5jO6QF96fGEF7k5mZOF5g9Jy/GkXeYF38lplclJubiG94feWEMgyS
odzM8XJJ4xo63g33SNdgkzlaSqEIciLSxkoq0n+raXvJtIlGRRmvQtHIROErYTgTeXqQKYnnCD+S
/xuOWFwIqjthq354kupA/yq4XM4q3aJHDxtRtLfqmDYjrp6OW3z5pB0RBeG0IJ7ve8dMrIseaoo+
0lCYDP8zIZkrIGHNdkPE0T/bkW+vT994hLNcXoLo5KJWvv16Peu1ZTnhF6wtgeKel4tRg0SHEj/U
KiC/BzDFkLvnWM1/QZx0pEigltfiq9gYAqSsSNwzRuWVT3m8+epdzN4LVhxSwyH8AETb6pPW6+9/
1floSkp+vAoMDSGMxucBsvrwWf5H+qMYvW7vlH3DX0lR34d/XQxGyZBCmb/LJw4V7B/mn+RrW/3t
30dz/v3Gun8PXxQQr62SYBsYKgaocazFo1K+U3BqUluxxMMR6d8Yo+czOQxEU8FvhxfIl8xtmhx2
6rHnRO2glIwpdxcy7WgDNxxn3IaTA7ouOC4cCHxxaTRS52+JCXpbnVp4mHESfE2IR2U0l9xeED99
i2YCoheOrzOCFM3LXufGR6vBLd90l3sqWyDiAr90deFXlxtIfNpbsSkvX2KWHBo7o5K4Pfa/vCSQ
di2HnDQbghyrJtKi2T/6dMkeKD80Xh+iTNFUG/DpUypLXpNk8d0zx1GOCK31t/4tLaBqCBkazjtl
u9XzSKw6pk782zV9KHprnMIgC2/GOKp1lDy2gVtYgLzX7Zti+Fi3o4uNSObfuFWx2hR7SVJoUUZ1
qnA8cG4xiCVVoj8MtfwcRlPSYlKXMvozairIYU3d8r39DTcjIacpTBxNgpF8usYXgOzvSqqJGIgD
ArQENkOmB8r8nYPlqy0mTQiO0vuJ2RcDk4/94c1GB3l38/scZyW7jk5Be2wsY3mzjA/5tO4i60EU
yqAd1YaYcAFpnxEg5CKmLzzicTwmrHqHqe4TLgxfrbtAvEMDNya+9Ge//uOHyp4gmA8kdmMWVogk
1urKQZSYo/hMWe4iF5GhuAUr7xOD0M+1ap7Bsqq0wwh+dYLCuUhIE1oT9rlPQON/KNKKcanbXI0V
6inf2dNDwaOt9PpFF52v1GkZPcS0aIKH/2Eqpv26W9lV/WrRxtBc8JN5lm8o3AvufVyq8+qxXoK4
3d37+kJSvlIkd1jvI9CZ/XQTJP+cxyH0b9TGZpChsujEvAiYp1p/cV6SziVymUgFYOi0zsaHFPJS
Hh2eaY04PYLZqp/KYfEkMhWuZ7+/T14y/pbVAh/ydGn69DZWFLrhM5Dl2422vrR3uAs3QgBdwjC6
A3e0kzl4qZZ/CQz45yh8bi/8PNS76yqhzg9wGnW2NTxYL9Jif163fq/7PznXPdR1DvrZPoBrB0ZN
TWwzA0qUDhzv0b7ZeU9yMgB4N5/IXrdeyjfanIq/MCGVBtw5nKfPLoRSnugxFcd8xB2yga6OXZ+u
eoMI0bituWXqI3/qBKtARVo7Y2o3jDFCSZyFlLIQDrg4tM7iCampwfGu6f07sLWV3OSRz7GOw78M
UFZaRAuBCS2uM8/KwagSxw2qOANO6DUiQ0vss1UNM+rtOwTd6tq9i8BnCmfrN1zpwQQNk9s9nqR2
2gGm0BoI1jA7a6+is1TA9hNGwxwH/kM6nh7DWZCyCaqAyOhdfe9M9nWIj7wAt6YLwuRwRIU3m13e
J4VnPXld0G5B7DBXi/ILYKhHknBhcQR6BiGG4XDQXNSBIc+0nJhRjLiKR++CSu7tNnANKiVsDEK0
Fph/hdgPDMej2weMkJVfYfAV9N25wBh+0ReoZWb5AtDWoPtsPRw1lwsTrqYb14oW9V+DzS1ooPCo
aJarg8w3Pr8txAWg409ALS5BAx0nf0B5+7wPRNtJH5esiHZYemoZGe10dUfY6hsPafY6aSkg6p6A
9NH9US1me11RcwaqLZoDs7blEL2wnFO3ekGGFihBSBufFn6KIsxXYiIDhGZpXxCx7lT4rN97xTXZ
Ebh4l9sC/hqCbWmV3dvJI3i2v2Ui/bp4+NFRVZSsQYh/oWc+6aPJiqUwX4MslEUtmSsGMfSQsJ9H
Ul/oNh6IkXgf1g5C7bgazzMx/frQ6loiJO9EjxZGLtSpYYCwyQBufU9m02ln7FOYhxxK0r6zAL3Z
FjH4Grprnkiqo8mN4Pb1UtvIpHHP9cyBLK9VEd7LkfNaGxLAFJYijgZQdTmHOW0qpZgaXkuTa7kN
BWEfnFVg4e62zk9d7ZJyzgEIgVfcV1/hYH3d6bAzs672SgMnHe7WQNamcZ5kvg8jV8CmKbVMGgQ/
IuPnu/qQqyFnPIX2H0NrJ3qb0AKXPOmYydRWazOD9JKetvk40i2HNAP46JOM/0ynsvlwZ9vScR3j
axkKOSXlBNiFiTQ2oJO/jyEYIhvGBzbQdtgjuSeT9CusGOsRM3JRvTBTCzh8/kRaCoaG5tSOYE8C
3vH04EL34qVKtaM5cJDlB0y6u8VbWKuX0N3R87/dGY0rdsUcv3f2Gv+iIcHDag5zZ+f/ZDeUATsF
/Hk/M2x6gdMiSaDc9lWBqOSnQNFgkVD6Fki9B4HWRcOyiJRqjbm/2KWLeVvVRsWFaRk6MKzi0mO4
evVDdvJwKYhuscBZpl55lNNKp5Wg4esfDDcnOxgHdsxk6fHLhQ94MwWh8BaYtU8wuKMUqZZChbyx
FcDp/Twih6fLCT7eD45RyqSv496jJ+NKwoUSlnGxxDbAAnd23JKwfTjNlA8NSWVUB8/79K6HqOo5
fus5Cj6HtIvSGif6Mt6SCBIyeOHxwlM1sKg30j2UOXpeObYcmZw27u6KTuXMAvz7V6eSkGryBlrB
8fTeNn6GqT8be69m39FCzFt0nokmU+6pAV5VimkfHC0Gmak0E74431Cc71m6du15LTdJsVeoYa01
WVL3cNs1+F6tvHmSlbSiVGJYnTo3TEGoj2h8UxinqYvo33Ztv85r+N5Zv3ETrDaUPX/edUAGeqch
GNsBHfWvWhoF1+I2vVC9DHrUaBTZnx5v0bsgOJgJENzHM+Rm03D7nEwuD7dVhM9k3oM8tCBO5IHo
RSoHFSn71Ubo9etWiXAS0KmqB446x6t8jE8P9wkAJI7ZnmixVfoH55e2MFaeCbUyb0Woso4DbNIl
9FFgC0EQlxg2ZhcMr+dMg2gwVVTC6xiAYkdZwUWLstqZxf6eHpBUsNk13soL9eBQvCW82KBYY7+Z
5aPaL0skjgFqHGn7x8JBPLBoCAol4MY4A8WUt0tZ+unufrz5eE7lKXvy0glHbNXkgxZvsf53kKeD
nSCnAWhwo/FrbkLsuCy4/yR5Fu6Vigu1eMULClKnx1hGFVpyd3TJmoIU7VpiJq5/SeW4KS+Sj6Se
QIbu+w/GploJ+o3BbVpoUXzSbHwhkWEBzMyd4MSebhwzsGTR01YbxMF+6fXnBewhKC3Khvu0rKwI
WDr3f/ZgNVHR8WHwQLIn+SURLPc67cXaOYDkwD8IhJQFgKF7551M9NuU1vOTYatrw77lC4djhDME
8uKgH52z2sKlifE9CZzl8/bLK6HJ2TIfa0GJDJ/brGXwANjfdVFsEd8pwUwLULQf+rCj/F8gLK5q
4lbsdDC6HSOPUlDtBoYLwwt/Sajbp7hhTGQZwhSx+kv1SQoo3dKKePAZZ7gR6HEbwWJ8F9H357rG
Yy5Xxhpf8QYQDnm8Dc5UpPXyhlrPPpMBow/1Wipn4Okcc9nvt5BjEuY5D/kFaACqYk0OoIu2wcxo
/vp5wRbFRQeaP9Kn/3L7Ku+amm/38MzbdLVuAgehOZycEKT0lwaKQerjuL3lGrpkuMh5wAkE01VL
Okf+hY3i2sNm7hppoMrB8Kdt3cVyifsdFDVFCKMj+CKWLi4+fo81yHni/zpHuWviwm4D3dn0Hc1D
gHASLlXeO3a+rIF/IbI7FllKX9xn64wT0hdMlykZBwjSo3/xFit3fZeyqrS9sZqAJI+ELgmbFQRj
J+/BfqNa7adgrc4B3BapYrHijVK4yyzg8F2xhkXC6W+uiysvlViDCiiJW3FI6gwJZIpk8bnSYp3C
IDgPp4aJQCplw3k7abHFFihUvAhplni8TR2hwg/IjcC5pgIKklWVyNQBKn054Nlz5+3JvnSFuUJq
VLJ7QRgp/Ya0N5wgYdJp8vbcH8XedulqoHPdDDP4fjeBsesl0WItgGAQtxzrNAHBDjAiUNxtPjTD
TJtv0NNoe9mL0Y8gi1/XkuOuVSIthH+7ycehoCnrBijpGgrcA3/BBWZk7wRb6YHLOCMrqDYFRiYA
y3WxFwgPHBr+ctKZtVkjMrRwO55Lreode+vWj0rSVGG06Q6+XEFyBcXXNoQOoMF05qFCv4KqWElO
YLztR1pGCP+SnZy56BV1D6jj4K0gnWz7Nbxz+faQ5XPloEYPLkYNmE6VAs3eWstyBxfCmeCF1m6C
7Bkmdh98Kr9GlOtm8BqleqAGza/yLCx5YRmtTqfwQkOgyKdJtkmUELvgziCAQBnrTO4n4cvIOKci
DsCleVROxRyNps7pwu+bEr+zoW0v/Uhaisd/K6CXrWVxCPVKmfO2x/gK8lyo73LueYslrnCCDL0B
aAnViYpp//meb0/CMOAEa9fmMsOpBYOoawiUOTXhHZGFtWgY/SDHVbCoETXK09TynmdRP3J8dGl8
MjoibvFRtYAJKHy01GhFHWZ2ZXqhK60FGy8qktz8rqGIbsKcf6Wjjw3uyHpFtejF5B99PR0/LdgX
5byi2RJCTkpgwDzNdb13ho7Y3+otfttYshSnGZfv2hRLMI/0Aum+fdkSnaB9uOR2pM9uNGUpmFCG
T1qpMNVFqe8vRQNZSitgqG8FeQXrZgOtz7t2+EW74Ts3Kdvp6byF18wU5kw9BB39QkTM31iK1PK7
fdMFjjqG/v1xEuNfZVUpEOvJqD/m6kXk/iquXqSsTEGvc5gAHxWhSzl4ox1R5B7ktR384HXqnKZn
X6PMH0Cg2N7HcNnbtyYSx8Q9LVBCxhmWm670YraN+Q9hdZqo5X09h5nAnNGTfaDl+BMRyoVi+zPz
uCWgkJH/ypM9yoWswo70/vIOlsiEuVBW5svqimY3IpafI6tLqbSuUPrr7VODqnSgIe6s2uZVPGm8
wViQZEGR5f0HGNtpF45PDg84RTkCy8gE1dkIpifMzp56fCFz8+qbEspn0501g5qjQVJQHGv8MrPQ
E58v1eLNCe7JokAF9nWLd9St13WIE6C5nbmS924Xi4DAGKRopEInJUu8dR+C/YqSKVOwGS1pbU63
9mZxeuPA+3jTRe+VBNhFuwTgGPAaH1H4gslC7ZqMQcwaurv9gbmn4B/NC0NDwZ2CvGRp2ymldDIo
J+iwVtj39D6CCo5pLQJCJ2gBP/WqKPLLe4J9W5mnFGNfHRywJCJ8jAZCXMQjf5uq6R1T76vyzVzZ
kmGDpL9J8QPs0fZfJdTaSBdrmkps2WlpvyinCjFjl37mvK8IlIRYdba7z54NohfCfR/jf8mETJJ+
8B6XxgMrvALlKfx2r6IGmc0cjRcvuNXa02+myHdQFnvG7uWeK3b8FRPvDdgrRh+9UGfhPJB+uaGs
VPoOUQcYkWjGG3lOoNRXAj/gdZPCcStyX2GJjcejD4iQz5f10yoTx3D/nuUEhyPSqOepJGSo/3J0
rIL/FcI0+LrGe0tC/ebhA23RdeqDpORPLj9i6MQDUErsZiTbCllvVmaeq8k5jwIj6Kf7zV06eeGC
rZVAQsJDCU6sLmsRt/AYwuJmBQoy4ia0Rj3WPxEhkikfmQ9NEij/MfNWPVzG4XNeEvI/3iVjbdSk
AaPwWPHjux85DMP14phVOQkM31HWN/K5h3QgD/Otw7EUgY8RT6vsjwFaC7rn0HjnwG+39wg2LDzg
Gn5Woe0Zh+ABedulPK+HemWZr8T6sJcPqPO+xuCeg/TyyraW8PWzVNNF3eFigT7ZAJoa/sktG0tK
Sx2iwfSfbQe2+vbWcDhkr07jo926kEVnS4NTAYA/x/rdGS3gcKrNQmWZC7bQxqCzd0lhIBsECX4U
t/cQZDl2ukyc2udM8Q1Em0hILkii5tjWY+HmIPbMNynvXGSQ+RusQ94tObskKaI040G0jHNsNBTv
yp8w1zOQAodWK0xxnUSk8+vTbxJx4voLX1fRRWzulV6t9tm5LDTOWbVyXP1eZDKSt5wemhdF1dW8
FofcqEMWpl0FUJxs5oAukm8/L6Xoz0PuxVSusltBGyZlPPzT76hWcLnElHh2xCyczfOcbXSrfg4I
M8zv9Rbi/XGuBCIR2CcS6i+MmsOPWCoj5IKAAbIp8iuPmr/G4uG7ETuVBaTbky4nmzAXGBx0LrZo
xpr52zMyfNDh0KpoycffElPrvT4qg7s26B5WACD8/WXpXaRkTJbia0K2z2ZEM+r5ol4XqUWaOHSc
SFNEACpG4p+Hd8J8Zr17WqwMOAIM0BoL7Bdh4Zmv598LXGGIpX1WrkL3l/wK2HbxKWbVDmYwYatU
GqmDW2zyghP3zSFkSYVXAIvHiSvwPfqgdjQNSv9BPQl0b55Ryc9HJ5yucrmmW6X0S3jZpEr1O5SE
Id6UZkKpEwSH1Vaojj0mW2bmNRSuxzJNsmZG5U+bKmLyfumf714L/DZgIqscHoew3AkbC8+DRQ1Q
fA4Pd/KIdE8yATapKfxZ6YK5hQR9FN41NYqGVhbrRZK6uYnXHK0IKJkLrfog9uv/0hnx3YxSaQdp
CKx9tH7j+kO9ss3F38VSBbWJogsr3okniI52r2zQCLWP0nG+kkiUGjoQGZPLMsUD9C4zM+fLrJ5p
Gn34IADwzKZpTIItlrYLDfWlUT5wjPaKqkIJIj1c70AL4UMiYA43K0unQGDkF6qzNqKPwBUKzbVV
wFr/+VpM2pNsySuy939uBqM461ZUjgQj4qBcNESdkaiIitWf4Ln2sRe7o6iFO3NmrRZ+PDKwFYac
9V5TSCjUro/ygjN6E2Nt952ow2X+BGI6QZHnjes3KGgXHdMngKte1lqg8/lr0kGpadvXkja8C4bi
fyyz7oT8gto7F5jwFtfF1j6uKwVfbsWbA3czRb4it1osScjs/EsQEXgbQhPkj2SO7D8ozITUiH20
UxiNA9v8xHJZqg5PCynM3Z9vYQb0iIp5VFr7fwMp1DCH85MVRAkzQ5lR+WRyXXUbntmUQpALgNjY
SWf/XdFUnCL55HJCyyS2nN+/CazSLej9H7PBsPKB8TBeoKKNnXmcuQgzA5IWDq1S7DreDRSkQnVO
LJY6KgG/MPlLCAcETvEfOQFzRS0NhIulYVOItznM+0FMwPzINBsstTwKhO+Wwd5KMIwxAaY7nPV1
NcERlPOM7Pq6Hc1kIGkktscxHu9WXIl5hUMI6UivA88kV4NiJ+jC8jydKOfUpGLdi0p2s0KLknMh
N8SHjTLXvN8BpSxugEbuiMXPyKn208bNcInakxECxYEkeuLrWsWUjqA4g9XTuzPkkQTNvNePenau
uyq8b8DLErZWvuh/d0RVcLKJxkYGf+82ph5z9FvSmOKgL9MjGr1FKk8p/pxzboeDxPJLdN/eVLqq
1UX4HV6mnu2UYJWjHy3oebK1bMRuc9So7zPJM/fw+qoVc+zEBUMublGPcHWZXVMBVJp48FIGNtK+
ASDDC1POUas1fZs/fqOX+0LxPyLoc3agALwTLyhlvGeR3Yu3hsuotan1MjhUJKGImnK+VbuFA1mo
pGYRVvoUKzxQ14DJ+xNmBwnVy/5tiS7DKemPl9Ry1hjuL8HIaMfraZ9vdKZZrDPjBIyk8UcCtuTg
N3eZ9rwzuPjUMeavgDl6HyASkru81X63ZKZh3Kt9+x5I503OPLBz+TA0sVbSxlL3VC7UnpI1Hy7F
6Lp+q7SJ8BRH6isrsI7zw97XYDNmJlWHZ7OWkqDXev41VQdrqWgYU73vKID/IX3UKWBAMZp6NSbM
u0QNiLVHod7TGs6pEqmQ6l900xB4tfhdLW1eaSXezl3ANUhyf4JZiwVQfGh3zAyUOXMd+/IIdYq/
aXzHEpx4vHeXGqaIYlxv0yMJCwLGJ3z6gv5YWMAPlrR4E8Hl42Wf8Ci7QKVz+558cGap2e4zmBDD
rDblBCfhNg0cBY8TYUywdF2o/7+5R9nBzb9G8T0o6X+Fjk5x5H7uTT57XUUQpSIyaxBGuS1sBoOq
2WEzzsXiR0Hhl3MI0OwhKSMw4eGA5yEaK9HiOA6jX0lHNnNzQtaTpwc8DWj5ig20N99tL+8VItKR
SG+N0VjXxce6ydYsoFAy99bBW4+zt/86w4bWZWS4aMbY/bTy4/YhcpPuBEPL878U89PLQl+/VU5x
dkMmF6U8+MkhyYqTGIRzNGrEoPtMPjjcZxuCdmwrnLVWfTBpWoDuwrnFpTdfx6BgfMg3fi47ZKZN
fC2j/PEsxtx52fxknFEGQv/oaf9UdKVLZWjdeuNWZCMyuS+9hSvrmFOF9/+uZLD1K6cKNp7eQhjz
S54EQnQw71LsXatc/yy3mOqHEI3nbVRR3PNwpVCy+XlL5+KhtiH/6Wz0AtL2a/2V+iEEVniMZO7t
m3/HG4Oj4hG1t6wiNKRv5D8iNJymtfPxVcJc++nyXs+MP5OHtrL3EBKg/+sZzF8eYqKTHn5vF9jg
HQEDXkldUq9zlPQIMcqdAB90ZUiXh2lYTrw6ErdaLnpgSFF6S58O7Pnnia88WwX+QgjEpR5Q5W5v
moLvrL5kcuUJb2MZXL+eUrKE0zl0SLDitgImPhpfgZ+BOpiHPH+2t73p9TWFc1qo7fnW/XGhPHpV
QduvW+PbY0Xf/WTxG/Nj8jourYR1+Gy5UxGxETdkgSknwluSe6oMqMT63u6zAvDaQjgSJlU0gdFH
bocmJ1PCKqCkFasrSK5DTmk7lW35AKKFETFW5xhlSW1YYo+vaR2BsqUM9eL0z1yFFXLqvCUWLHIt
3oW+EBXc5Bu2G2FLezAJjR/KNTXyQh9uZXilqUAjx1xZPx41xl5ol6ofioNzwqbSP25R5R297G8U
P81JQoBvbCIxuRVh8AIbv2BqS6ZnJ/Fcf87ZDg/QK6e0rM4OgbFtj4GLewWhVSzdRALJ/dsEc6WH
basZO4XZdb3TINViHzuk9ZgIDAjtVDtUATQtoHWqGnDqMLR9VMl2DW0rHg0rRppA8iP6SoqDaNYq
Aub5v0G6moziQcDuxs3q4TJtVHXN2qhwH8T6qPeNbvFSmM/WMc+ad/MSGFellawSLTFb77lvfFzD
bXWIwi0v2qjmlyRR6doDe0tVEyZF7r92MMCAECLOTMnIy/LEgRx5R0TH7fkO1Fwyr5DXdd+uI/x4
p/h8MMFJee6Oh5k3ZlCCK1VwIDeCo3RmMWMnry8yE8KvSeCxsusueSsqfIZ6robs5aVs0UcY65N6
PeOvc8SYdhNsCjoGHNYajQqeu1DUC50fMoi1RwghmKUefb/7U8jsLFpfbkPugG+IP8NaFwS8yRnr
v1n3MCjli4tLNhxxza22c4/jc1/bsz59i1qgUlOdypCOQ1fO2jWtsUdXwARqT1YxsO8CEzDiSo1s
wjQMizHTSv4yV4z30C7WyaF+VNAmOUXTkg/KfJe2A2vLw1wMBxNk6M3wvXGm7pEiv05aHue02dsU
HeH5XdnI/Gx49bC8IxtjTRMQXZDMSTAYii0J0AQL7NGmutr0u/pB6umSrfUVMI8kqdCgxfSbtrYo
9/Fh1g91iPzks4jeyi5FsubTBLiv2+CfcaYch3toVjL70domxH9iAqfWVMiq5FUTa4sUk4Y8iVm3
+oM8TzwiRPQ/O1WbirU22pRywkeNCaYpg/5YfwNy8EZSf/HeTy+Edz1sk29B0eFOwFcP+u1lQN7Y
BFi2cjV2p9e9PmkAf5hQQhX2xLP2OmouHecdH15G3ysrl5UQDUwdUH1V55+PnpIQvA+dqNQG9OWf
/qxhMCVBwegw7q8KJqICPckwqpSpeHUTIOOdLWQs+sxgL5GiFLgwU42RhPDktErY5MvTSZSnigBp
5xZEH3ThI9U7zMHkwrfGzh8vaa5xcV2vBzn+JHl/kpEwLFNUb3LprCG1HFyDZ4j2Tr6I0bOhX+6T
dtSD550XyXNi1hp69CZf1jeVFmjdkvktbagvZRg1fkHfKM3mzaMvXl7MjDzVGp3iFJJZFWf6qMok
BSKe0MaDql4twoRWx9cjhcn7+eJEZcMXCA4NThviUNhwn00ZIVHa3GVS5tm50vbZxLWb4uLD7flr
rfE7PO0EsEpribrCmdaUb4h31SdIQQbih2qWKwRn4urbPbmxVTFQQaQmL3SMzo3EUFmaCUaSqZyE
wbqlGESOS3d8xzT+GMF2I5/WexN04mmicwoVF1FQLIWltOwZhmIt7cIibbzk3DlLNfyLJGw0ZSmE
WvfD1OAKkHqaGwPiZXTwVvkDc/0iw0OqG6n57Gdgit8ebJ4T6i2fygo9HC5ymzivzQ5756TE9UMY
E9Yktl7kvrwD7WoShNnuq1l7FyGitmJ80/KROvVByfR2RfNHrLahaDPQeOYTF+u9rnSVeUP2X6NP
BnrJACam/aQD87wTHYo5Xj73uq9Mdp5EEvJikTxett/yQB4SQAX/1HvZcA5CQVtWUxxE5qqpk206
XW2ZUFQq0VHFkYUkj4qTDvGbi78YCBduY8vd9nbVv2KQmFrwJhEmtv6iUVEVc2sd+0WhdKJdvYHC
SUf/fnJxNIcvnH9KEs5KOfHKHp7rQAWANlLRUlbhKxru/0d5XMqZBFmbmvxE+a1SAszqbjJgW428
DbRtCXUbFCI0ZYL8ASwLSv/YfIMBFIg3LHyl8/CXt9rzCjDadn+wV4AdfGIifVBV3AbdwhBJW8C5
2ESUhjS0LoxqF+G8IX+/LNNHni9mEY+NVk99IeydkVpEdCc0llin47X00nr1Gfw98hAejzokKeVe
VPwKT5LNr3gg22FPacYitsKpoPRzVMheaXkm6utfo5ZSPTSQRstNDKFr1EBCA/57lAk69MOH0AZI
9ZLK92Ppkr244BbKCcisqrk09IuoonkmGeqvO3YiVWmwyzc4msqm7wQWTSKYuZ6B4FZ2ZvgFQzqm
Fu7oVV7O23E81yFGCVgwdnSrOQjfY9shm4a9gdGexOfPltEEx+RkyI9M2mdCSoexwybUYQ6i3cD6
RBuzVPFr1A+eXHF2x5dvnko5/IrJuW3Xq9DldygtOf1berdzcbORDVqCAaXBHkx9JwXz35Tl1sFt
Lqmy86jLaMfZLaZ34MpfTuYBJxx9ZVow8OL+m6dq7lkeXBjFBZn2J6AyGKGmXyo5RS57doU2EN6R
xGx2iWgpymrn1mgQOaXC1sPaRBUiN13OFiAhJH3HQT9PzPMzBxYM0AVHJtaGy16obHpdr2B3N2oS
fdspcbtnrOpKqhYNCivS65vhiCR5xCYBnRwJCEgPmVz3Fo5e2xtPTJFoLS5t4PfUO8MksTICrwnY
89LNDHbbgWc+WWqCCJvyKhD5ApXScSVjieTTx82Hlmk4U+K0zY33isBr8fUCG+nspF+JK/CtUI/x
yJufNFYYrybKbhInqPXwvY+MjdI+Ptoows2szmqd3BnB0v3U9cZt1YbGESoDLVsntNBrce8kTKV0
SSMqkZ5DwvWMR37JVggYfcyRnjXvAVPNhUjwaAOzftG0bJ+ENjX1/0PwIm0Hubia3VzyGt5XyOB0
IHUJx4+gvjCOCDuJ/W4zNCfEVeLCSWc1ayUnxYTwzYyZxuRpDDUVNK1vmPF5Cv6Io7kozEmgFScV
l9T0RB/Z1tImkYS9knnZ7u/540aKy7OZrC8/VS6f+qzJA+k5pmYmRthH7eBv7nYnJQiq8zaXLwgo
mu3nWNiFJA2sMXhoVY5YNkUzE7ItVeyvTiqVdixjWTK04HTdDIg7R0BjiQ30yepnSegbNyMjKK0D
GoszkxDhzOcd/rCYFB19On2KY3BZ9et10L9E1/ae0KktHBem1db17LkEISr1Qi5qymCj/W78pj7t
5RKDNEUzWrj0KNa5EZ2i1307Dz0IK68WbL+r9ahClT8XGuouOjmz0KEXab4cJ6KzVRzYaHInxnqK
58QmQsKgIkO/QHLHwBvvoPibMFN9IKoaiJQg4DtR9ymE8uaBkB8htKS5rarYuHGfLQJfty4aUY6C
G4uXR8+mvad3xLTIOgTsXEuxs0/nt1VDuPewtTXrGG7HBWUt74XheBlq6JjjlVsocc8MT2f6frhP
fL+GLz66TF1d1z0DoSzqICF2aPge8UDqjc2CivEaxc9Y0wyUNQu/2Q7kh+f/L+wWIYKatBroi8v8
mtb+u4/c4KGXv+jWmANMK/d8rwGaOPo2di66s+0f/cHUXPAkUz9MYG7jkAK+N5I4Khem5aegYKT1
RhZSpgen026SDDq5F8bLGU7iH30YucB5AwLzzbZH59bfHFbQ7Nb9VrBkuoWK3ss7T7I9G5MQMOXj
9ENuvq0mz/CtGbUQabUKSzjwVl6LZn6M672hJdr2lDAbJW7rL0p53Mx8p9Zr+nlhzcZXy1wf6TuC
noDVR1wpZb/QkVFrrQUwy6zOi1CDR0/RfmG0Ifps7qlU+7iFKRkvw1Njrlvfs4qZxyP36dDgsakq
cxgNq8m/dRjoBdyd9PEZ+SxzL/HsQ/yfDrMaqE32HA6QaYogbvgt0O+MYCy8z8B/gMxPB/6gveXT
t4AThbt+zamOSYD7jNo2t3b0R5Fus1k02dXQgNU1WHxm4qpEwrKP10yEJP5+qiRAckKkaZxL4lGO
KwOXqCxc2cWd5Y7GDsuYXJyoL/28HuIJx5Rmdy7zQ+qsq/dlEg4DX2mcIcbQhGdzAdfj1STi9qSu
nWtjzG1Qkv33+RUgEjlnJtp/7b25SkBCVNP46yJmiLqjDiGqxbLIjX6yiXNzuNy7hrWYNDJOfC5I
rBX0kZ4h28sBbSgm4VV5p+yZcq304WupDXGfYZjpVqxdeyqTU/H7g1TZ1M3hzn9GCw26HB+fXaoc
Dr3XmwYPM4il5OmlSWPBurl8omlUp8AuramooZKdBMO7fYeHUGHh2bVVmORA4CIWAeqYufrydcSC
PSK8X7/wV5GQ9lER6Zr5Jt9T7Ld36kUxFEVAn+z7bsIMOW2o5D8gVJJ6xyJJssNxnd4aX1EwRl+W
TvDFNwSUpDwO8WzEDFVGhkNn1tj3StdQQLqyldnInk77wdxntQr5mSHsxRO6c8SX67RZrQ+dwnSU
ojsCsG5fTEYwJzlZ3MhLdYh/pRVduZX2+k8jHjwJnGyphBQM7n7Pj9hWIKVA4RowDPBWGq7erBD5
H9NpTLv3WpK9gpzXqp4F3gf6+Caif9qFNO3rHCspU+t/sUw45zRpknjrcYppxzzcTYgsWY+55DBT
wutYuScMAv3jvnfczddn/gy3+aI3BqTLqX1OdwyEjGK1PxIABZ9HHCoRYxX4hSkWPBmd3MhaObhp
gyMX3yw83tqhgZyj+kMjZdoyZKjZpf06HLc9kZzKmYks0rdB6GV7JYzJuUDyHY6BATSSo8rjQIzE
rbQ3P8cPJDeevheAkOfe6PheQFFZzfubB7L/Cm+wrZyna5J4ML7MEX8L1pVjQF1w2Q1wmxhnAP2Y
J3+mK4MvXI8bmG/aPHBlWYAzRo4BwiLshvcjTzuVAMqCItIZHkf7XvSeEO8/yy880dLJ31e8QPCn
isFOBNKUceUQNkFApPmgiFH4VI4qiNtb+6dvBeDZRaUgUb6mUTVa3i7yHWt+Mf4upV/v6GQwLEHl
Sx7ZfUOgC8HFW9xjg/kIrtyDQDYh0gsdaM+ziEvWgm9o956PktNmy3ghBo1pkUvZEaVjRKsijWC0
cd6E2KVIwj3zSG3sjHQoRHyeUiOgkXSnwJQ7zJED4ajVEKgXJJdMHbYZsGoVQL8eNu7QExjaGXhk
EBu6VldtEyhK8/K/WxVnYwX2omvKtUXcCYB87OTcAVviOKRfqLEXWmTzJH6abf+zWEfJxUIdTS9m
StxUI2NVRiZU8zzr1ZRbv7BushDXgHeCKScePsRcbfe3tCvdw+8cg5Y4eT+M3LQaMKJ9D2cF7PMs
vA+W/zx1bBG2Bkjd7nbioZqrM51ZVCs0Vb3oYXvCHqAq9b9yRrRPnkhFv2KKvYtC3nwlaUAabHsW
WTj9g5KC4vKooC6GzbXNnigN6U+qbQAoq0L7FZRe6y0tG52TAbqEvUB+q28mzVLHI/M5YQE94AHC
yrAUgaF9RvI0ogg53xrFf2Bf1252d+CIuPp9ZwSAPlvaNgZ49XzZbweGYJL6kmHqIoqkQ47IEGuv
b2HvH/QhJZxRF2jrsKR7J0LjvW12SqLD5fBlFXINQVbejESnDTI5QLauLK8zTeU17cdmFyk76ziK
XhtRasuht0xZQI+gtEUDJnuzgb4L4KFrT4qiPkb9q6VZZMga6nbPkjqcT86xp+aDI7nlTxhZ9gfR
2cFdB9kKjecJt4v9HoRLegVP+JKUryJYfHiWbBwTeL+Pso8MeMrMqE0wt5EDUa0gtwP7igl8VbNG
4aO+GvfuCmGlBWdueIHX+vf6cc6qJ+4pd7kmlUTdb5MuNxcdEj085Z6kU+mftdre0mVoSZyZnvOr
N+M4+7gb+YLKkfVi9doi/mHWQV1GUyZ+X3RgoYrgo/l9fnXp/5EAxXVkq/y3xSXV5dgmG5ADEdf6
nZ6d7/5qwwGaKIZ+0evY67ApgeQjaBHcBpIW75kWL8oIhN/LkhyLW7gbFA0EkmwaIftxzXPbD+a3
zjR9fxPSvrFH1Zoh9qo7AoQbwBYT0IlqmWCxbxsYHxlYPkeTIK4QADQEFqgmgB6UIeh8X75dkAuq
+IOYm5iF0443tvHzpqa2PBZKvLwLgJQBab6Zs+xHBYoaShcNMxDY6PUxWwDlsF3POL6ltrtjMepZ
p17a7ftlHo/Bpn6VXLXq0ZGJzpQynrpVVm0Vkhy/26nG7cWYVSkpAOVxQQ9qWqq25Th/VrBMf3N9
IA2BURyhCqSHBvmYDP3WKeZjq/8my4Yjhot8eD2uJrKjYva6+E0KfJoAZ/tQkVM+TxHTySNhOrdw
dos1+zpwIhHoLhmxhOjBW+ayji8m0i1/sUKb2+Bjfta+8mR+KxC8QWSh9PCtW2pLvGLipZ3Wse48
HzLiTyWs5WTJB6fSYVHti0S8+SkhgkDLKqjTTbZp0A0GiAc2vF7QeIR42SMThsL955q2l9cR/QaK
vzydL0OYwA+ecaEKrvpr9ztuQ+El+JUzkGcxl6761OIS8rOOwmN+GVaDssOKX123Rh2Y7QjfrmYH
r174sQJksO4B5yeSYbEyGjhzvpl+di6td/tfAI9gmCcfWSrKeJNXFd8jaqM3ifGWqB/judVNzJ+8
3GIpBw6rPhjsr1u/akMHzvGny67Ke08LaDmrpYQ8ziSl5XHJn1O2m9pYfKHbTAv1qdk/UNRBSo0e
9XMWP+AtyglErz6iHBs89aI+IyopOmm1TTd2Zu2w8OR5d0Am4naMK4YeRB7LmLszWjcpAcqGLRSS
KUdxhYFN4T6pRbNJmuzimfZBD/J5/rX0gB6YVpfQxr8d+fASB3ufIjDWlRKKZH2ouV5OkHc0lnTL
Nwe/BJp5vU7MPaSkBPKspV7wANIO7H5exQyjfeCu/aVk8cnQ+X8vsaoZqNUfZq7Mzryi3b81E6CT
/AKw1/lMdGrHAu4sWWg2hTSPpcABFa1Mo6lTRXjQpTVFowrx3YG0dEJOunDPHIu3iNqsKt8/YlpW
kv1sGrwSR/nbjqrK0rgqIK9uhd+D69b1nvX1i8QqZOfexDmc/yv16vTuv8HUO1FeQCqq/+lJ7Nd2
FkjWJMbHEv/f4ZePR6a8hH/T+Rys50CexkV6cglA5OXIsElqyxBbcNQGKnLIEkIWsPL8W7YtueXE
LL8j4M6b2l9H7wBFmed5D3izw+baFfWSAVS1c8YEBtBajMF+f6rcrZQWlmxm/O1Hzo9OsgQI9e0n
gnK9unoIaz3I9Iu27YbVfNEQsvcOS7HJB8AEkJhovhSZ/VSCnQDibwWVMmKK378dvONz1WR95JbM
aKZ2mcbb6IUd5QS4NjFpqO/AO9efWWWTtCmTY0DaPXl+/8WDBT8bjJ5i4H+PjlKJ80zQkOei+jkP
SZ2C5p8HpkYBzQOy3hb0IXTeUndNfLaEI7bCI+zqf2ymIWYakcdb5FdgZN3pdvKD+6nq08l46xC3
5j0ojYYYRFw1D9ThKQMRaf8HMySPJ2MzvxAT8ZgkGVniGFWRZH/X3axjnlsgcDdLMQACWVuVASVq
CYZqg0Yhi6/8pNVPwkX1UI4BkoGUi5Tamoyz1Z9o8BXPKF9rOhkSTsDYKvJX5/SzP6Vdsv7mK7bh
cWU/YEkzfFVrbwN5xlDGfa9/OSuOM/AET4Qt4ioyyntZWpRTa/LjPMOR4jSp7RpA5cyVngNwPa9k
64rlmsKS5z0RyWWW7fT3KXQw1SRqI1EJBW9CgfTlLZVICnEBTx0dlp1XC22YHtX0BfH+RxE/Mr8+
3/IrDS2XQOHX8/Fcmyn3S463nGcYFYZwUcObe829IDmTjzFrgOSKVpWzI6mdBnxAVRdEx12Sxp3s
7tl/+hxqv61YO+8kzJHmv4MCQTduJT28W4wb9hbMVhL4NIk1bNqDKO6R1dUZ0mqQbrQbPpY5JZq5
EVRWsEV/4G1GwIp4+LzPJzE0QhOy4FiJINCK+rQSol5MvJb36nNbhyHCF80QBjBWBNcxS26BgFbC
JSUt2DyXOuZ9eBFuw17QfTvSDo+VT+aB240rXw9EqFnT0EE6G46eGnbupvKml098lDhBC2EvMMFL
N6TdSacXvXg/CVXWuJFl93CG5bMWINB6zwqYBYi5Sw6x41wshNbJHRzvTBkRJFAvAqVxc92LfEl8
teACpmX+G17As4h22+wZCG4LcLe6+/j2RiCDfQst7M34lmMyMzOWd0bj7acm36t0zsdchbXJkOiL
G2RK0In8S54SFmgk0RzxS8OD3uXIqj4zbavhU4nZcHyMniSfR0nZcdhpTKs9lmewna+xhDQNwgj4
EzLetcAGlTF5Hh3FT+utvxgGIvYfb4LCqJiYDctqrullAZcb9+wHcbBHCkkUWS+P3zKM1sLL9otX
mJ27qcEMWmaP3GwOHKn6Ad/o5dobn5y4f3sRmbGZWZnXHnQIJIEzONyiAPOq9vGaNJcvRkVQ1IdM
E1Bjs2WWtDmLzaN0yI7AJt4/bmU7hKdvMqG1HB8YqKL5lww5oZtjf3MX1XLM7NXcE3uE8U59ayh2
jLC293lG3I/vDFqyc7tVUaFJnxt1ouLfbvmRefkO6JJ33Z2souxja70sSl7CJfY8os+o3HVhd7m4
i0nfPiwPcXYDmWztqZU/Fsepa18Zh6zAOf1WLm49j/Y/hWhzLMe3St7H3ItsNlKlug94KLaI7c2d
/OOVVYSRuhgtde3FnNuIQs0YMRm2lY2NajTVC17Tu0HWG/Z+4uK+AB9wZhvv7T3uwN1ksxc5l0b0
dDq0h6Hc2oPglgnIHRCvvxQDl0yCOwCrK0Gw8R8nXN2xf5fOtI98ne/uyKACw1RfhogO+EdPvuJ6
tb/2r8XrsjPP7dam6lNjMcrleOIsOfpMnqwwBem0wehBVkARCgQ5dwCz9D+dOKr82CvPANw9e7y/
6vg3XUdSot/Y2IRkaRFzwKmXA5ECHSQJQVlSiJJc7qfkbJ4xQFZOxbn+7iq0HRm+JGKXQCYXInFp
UIzItHWVf96fYlj+j73353KZA6/hCV7DT0IhRVmwRxmDi+m6yRta9R8XcphmC4xlOYoHmtcW8shv
pNa5r7lL+evqvWLdfDxNy9J92Ju6PtQeza6dSgLCy38MYk8PgIOeE6n5KDkYRkAg6xUaCD3y2FsP
Xa2uqaztyvof0kfWXqWzotFWerQbLli+D9c4B2dPl3QoyOJ2/fLoHhIOL8f/odWcLaFPcudk3S8r
rO/ykCQ5ba5Y0ftJ/sgtPqXS/1RcuenEkCuxyjxhTTqLFQgV9sKKt40vAmJ6lK4Pd11LvSkvlCY4
/CYGNAuBmHemPM1TPKT83EWwBo8dMYtxY2fuTeIl1Z7BFBUHxU7BZCjNZEIAQb9bVbVAaTOn+gqL
iLQecr6UVZegESu0jd/oDnsMxtDGgkorX2iCfoWXmJjdqRbfeoHWmcvDQAfuDTmtyE0MQmwEDwz7
3aj2sLtgpV9gxm7Z7FfQDgpRwSb5f8baQSfmDC7HyTImC6Qy2dmZ2qdYXZGPM4p24NMkuMn2ewWd
zV3kGeWhLWrBKH9Wl7ZwgtXPfeNfy8eH0kR6ADktjrhCCWv9Yv+bIVwjUAOVurdGMqlB5V9wwewV
cefedFg14XAOIEwRjHtW84EP2QU4kRuTzTBnQWc/JpD+i96VSAWuFnItloXhEWV5BKdMs4C+e67C
zwIJLbDmq+lbJb+/WNFt3vPvroyYQnPqe00In8RexdwZ5spGc9coZjtKgcFXS3EnEuddh/RGvuFM
QNKnU7ZYwERZu+1sL+E3tQYP5COeAme3NP7sCj5Iwc0uD9Kx/QL3CcCIpiydMuH5uFGpKmUXoek6
7oZE5yAInDrX5rLe7JAwX+zXO+B/fRXgXR5+ml/0/Hq5pmO04NmMQoii+sK4sFiGXqdaRLVgAFmF
Wd7mP0uPcNXjMFpjMJgiLYqmD4yQqAde9fnu5njNKd1ILv3Hm7I5hjGEXL5RTsOrpdPMb6wsQpIU
n+ww5cHnKHeYH3TxYpoCVU7AHtV3+Tz28DOHB+tYy4EVky2br6mM97v1FPi5yoEN3lmPLGI+fXQL
sksvxuzhE1J4hhfBQPQpD6WpJI8QQpmVr10iYoCv9L/rvkOjVtMxs6cJZw2MWlmYPGCM7Ayw7Uwr
SINfQssWcx46f2p+BTLB5dN+YIysBlYKo3wXPAOWskSU1YYTrp24fJEDxLt4wj/SvSdVHnXYedvH
+gDbzELP7nKnj0IqZHIhGGTcEZrpsAE+RH/Nv4Or7EaGhIbv6gW4XO1OPBiLseJ7ZKL3SggsvRqB
5CUJAZTW4nRLlkjV/zRBJfdpnWz2kkYKqCZd/Jgv6UfXu+zwYJTjlQn6t6jCCSYxXjPlbPKzBw7D
vafHiZspxbIdxF/H0umCpOW2PpZrv4/zDPEVcCO7oQEVFp67mGAj0x3Qu/f8HIYNWsFv87DQA391
vMAV566XFvqXolXSPNeWJWU6U5RG4nmnen0mzyWegxbGjDE1GtxxUbgWwD5rAWM04r0yfd3NfAQ3
lIwWYpMMBKuIQmUvximAG/+zn6xjqGXlTcEzBjR/dp+w114Ldk+NWkWZjyp9nByh13rflY/CNPy/
3qc77XIRcTu4Fv/nwDs+1a2hDHIDd46PcOLIj6Mad+hBvZf8D1+O0C0Ve32oye4ncr55DdhvhlZx
iTUqQNtOSARBtNGcIKiNTFB0UN13dwK1olC9ml7kt1guemsZeO9jK5j61AyPBwN0v7rrzg7Et9DF
aYbFcRnOcKNd2xMdHVx3CyulVPGsi3rCHwXqUppYv9sQ1lg8y6co3zVyU83DrqMtSrQdG1uG6WCM
FpuVhQC0gap4SdVpiCFtQY3cmgXHXPO8kWbgFml50ASvWbA4Cl4q4aEtUmv0yxlR6RLGKmsVwrSw
rY8YnkmSlQnAyR5nalnBcr5KR0o5faGIBr04nP492Jd5uaeXufhV5yfXduI811dRwjalNJFLCRKK
P4FDzLZWd/vtpyOgEIkTMZh46g/kFWA6OkQPp8ZZeJvvKBN5piZlEpuz9t0IKWDcSE7D1RZjMkXn
9d4H8EvSlU2ysU+rmFEPREZGvRnwiB5taV4ZrzdSJaLlFU1mmZK4JtcC0FdDiuN7Up8Sg6Ydqmgp
aE2kDOrsUYbY8KZ/hS4EWXR0JbEdQY4nX3J8DY7mRD0GHxms7UudojMymsitrwDZRzDhavZw72g3
KQnEuYpLUdGzzITEx7oiQybHdcyw4UAHwoh285RtYgbCFNt5uZa1HUGZeW9fqByjPL+yBXDV/o6O
oxN5G5UrdS5OFRemyl4ncL1XS0CMH1B51lsif+C4saUhfalOysCbPSj4a77HZutaDvapeejM0zrq
riAPKpEz8jvgyYshq4TexohxHqXLLh3Wq8I0ia4YwhI+8tNY+NoDdhX3JbmwTgd6eB15ttw1BUQI
607NjlgiZPLqPw2VUcOpksmP+lKxsogU4C8EtYereUb/SRibFhAIWHFiXO+jY6P8y+bqAakbNIDf
po+breerKkVb7Z1CWYeEmrUCeP7CXQy85oZr+DRalj2lJppEwSxhaKAiK+V2oi4oqt7R5OEDZZdn
w+uMazbLiInmDakTohfWBptjHVCb+Xxp/pCZCHF1MHL3fFoG+5U6U6q4gZoUaMi/h2h2s2y8IWzr
+2w3nTyaUALkBpY5l8e7CyFQvfawI04JzESJWk7I0+ytvlaf4IzET2RJh69Ys6AzygneVumgPHCz
gWD7ZkWG0oNSEPVhfcknOqfId+EAQpYFbjZrcTeBJvYiBFg4EcuGHWQLp2lFCLcYwkk0G5aowMdB
/8FuS04MH1HOwnU6es3Ih2XIhZStc0Hg5YnzV09w2goteLRT7VEqw1Qwkoj+S2DWkxxhxYXo2XDi
zUHol2wSMsbTt41Se83CRpQ89BPGqN696h43bxM8BJOEmFbcvegCTgcyD/DxnbeqAwD6f8RmkLLe
bFuWRsekKNee6PvBR2ep/mNVoxXzCP6VHELYxD9oobopoBwqUJAbIKSQfJ4KZKobBDy/fWbfKFFY
pfIpEMlNJhjZUulQoCCL7MClKcCJVZt/3X/T/9GTwP+itOGtrNtO22G5jl2z/14CWhB5xId6CBFZ
FtjsDtQiT1R3j3WoAGKfIRtIwPJdojQoFgEo+TyfLWOYHq9gyD36CxjLwVD3vJ2F1h5VKlxhZPiw
rJnEIKCJTEh0fLeLRzDkuneaA/f8Y+NPDdP08BMr//joxLfkDdSLBcNvTLAYQdRJpie9DwUn23QX
k4s02CFB/jLYfxrOFX7+SWJ/iQa57ZbIKVO83MBytBXh2gVn7mLLe1GND/mWFgHlAvpGZNMk/dzG
Hvx3QhYY0oASrka+AvlMt+xcQ025/vB2wezvi0uHj+YNc2qkiNATHo0iRDWoDi8c0ABas46OeYuY
lJ6hfanW87J+XnVZ0zUzMRWjrKhhFiXSOB52vm0Qy540NrgH73Ybh52g9buI5mKAgQjxxN2MCydO
SGYWvxD9I/hCEo3npDyLyYDAKVjqOsUnZ5xfFtgDJQhJkjaMmYg5pV1QEg91SCZc2BjrORI7wRXH
ECu4OhXOPCWO6In7Hl47NFe8uGiYrezL54n+inE7vxxquNdnYYol0TlR+ivkGH9k+aZqa6KLG3QM
G/X7VJwFLweCI0GE0HFkkRCnRQJF2K6F0kCGy7w8prmRGm9mKMaNj5z9DRemBWv5K+9djjXSgG3g
1Y0oZ53iXw4nOnxba0vDP2jRf9sciDi9kfG+r8Q/sR1L4UMYCnhpMQOBGAG4m4KpszNEH/UE3vLr
tj8Gs77J/R+foKJ7etfrb453d0JIeKQEqO/w2+old8Tq6sUFHBk0/tyCGZWs2AmUONLoKKQvJ5PY
4JpMTvjTbEq/b5G4vd7zRVKqf+7KRpfG+zbQ3vBYJYMMK/Um9jbycp9EUXmMEXoHvRR3zTHOcdjz
8IDqalY7y0Dt+2ageMF1bSinaWY+uxitCBwYizCbsCKXD77cfji2mcNJTfKncjpSQJvtEDYXXXAH
6hbcFeLG+bTqlJJD31V7d2B1O6A/Hi+v8IPrImgP7pNN4nbVf96XvmatOZFVrQWZ181+4U3g5mnr
0rycNK92Kf3PMQ8pmSNRLVyshm+aNHS9QXPPMyMEBvV7E30epjiqO7KPWXsSjYPpN4ZWO/A51qbU
KKVL50xGZXrjynziOzfBcFT8SIhDP73b2S9wLiYrGtT3wWNyrw/vFP7AcZnffSl6LapEcf2g82Kz
c51/VYLkjajo4Ikwmqs15troCARC0j7WKTXXZDKQ8nJFhhWc/JKlCYmJWfga2E6djUAvbUCtDBe2
zPJpb5njZqxgL/ZDaSqja4KS4BFdk7918kWcf4eMF9xzpyBjtDGA7Uq1218GxzEgnX+dav7aDY+E
E8EE5TYdC7hFEiHLnBsVI4oPf7yG4CJfvNo5CM8uzmnoDPddnlCM+FsHrUUi5CR5jnPP9ff8F7Pi
KCQMZJhSrHKrgBZSLQv5Y8bEGEn2t9Qp8XGD9XiyMJc7ydsYDS+u8FzzFaarqb3mAkyNguXwjkcL
+mW1FxefXZnrCj+Oj8MDRacgB3Zsq8cEgqtBky5eGHPcZsJDk4D+E54ByM+vUnGhWjCQEQMzGBtG
cD2egf7sKZO3N3zqv5dn7Ruk9uSknrArkL/HPZNyer6zlICsRrEp/keL+ygC1UeBz15Pg4zf4GO9
OBPtUkcJp47IGJpHbPX9HbvPL9iWoV4SHwQI5EMggirjewEFKclg1r/LeycRSrvBkDujitf+FEVW
xColDxlrrToF1jqaITnNyXMker7da74fM7LDA2zLmeZH5YgPx1SLFXgqS14rmBG2ISgpxtoMiZAk
QCB2yTFE4IVCzPBwSsfG9iHUDVFEIbuZ1myocWz6fIAXTVl5E3+3FXNBIxHn/E64BuGIenmupPja
nXuPaxcVpIt+UAP4NykRyQOYWQ2SIyYoWwWSCX1U7Y19dQ+ANDjnkQsZBbpr66B09YWhT7wXkfx/
jmjnLNFpBDkhUPWCtKZZUbtAN2KjB4LP/pnmf5M3ihn6MXQbLoIWez2nRT2K0XhllpUwhsz4w493
myiUKkkzpcZCbiuXjK0L+YMBgholcAU+SqYIzVUZHqsTB97IGCTx35z4EqnOcrj9Bqm7wISvfl6Y
dgbtLaT/STkMQe/lGHipuC6fm3WJw2kg9+VJfGarH78AxMVc9Ud62zyZrbEZ5aV+qyLQMnRukfuP
QnvWyWr/sugbJujU25n4w3kAKGnwKz5WL238vK0io4lVm9yb65YToxj7YHiqNdljfR6fqavKv3xo
Pna5dFdX5fd2VBPa/kJZuE4Q/Vyt0eyfqkxqhIeoi1uOo6Gay+miHTBGNSP7foqxgyC/yvXvts6D
IbcBs7b5IR9e1aCLgJO6UoOwGLLGG/uXwcQ3WMiGLkNZcZh2ZqJUKytydunEKQzVVG14F39kUlCU
x13vFM6wHybgnSr5gec+FfeatPJUjWhXBcOEfRCVAR1qBb8pd7/K/qv38nTQYk5CcNH2RxlPcZHb
QcN5f8FpwP0j+K8189ub8SSY3qtTvtY9odl2gzqW/nZ3zJeq38LgMO33tzpr4iy0O29JFzxZL8Rj
6e1JN/+EVXPW6x11FsQpXkM1DMPgHkj2VaN40JjRnA63OOVPP5r8K4roAjRSUomEIjubzMzdwxJO
EN3Z95jbiHb2mq2+z7CIkuS5b52I1OybNUJJQRMenmL5rn8xGoS0gqGlY1Z1G9D8Akn7T7axmLnN
JcvO46FQES2Rsmf5vszmmW7t3Qqn381JMZfVgRfs1Dh1EpD+FzEHzVblzaH8fbO+aAce1BS/Nme5
7udTdCfX6oG26YG5Re5350sm8xAofNm35+vRb4KvTIWyQCAJB5Jcf5W2XLn+GmFWZDp3ebwUS2F2
o8S3PHSDzpvnPXJKYBc9WM+IS+aooVfDQSQH3cvVxBIMcw6KYoODN2hjNbTIzJajr1RUTNAVW8A5
DIpqoD/ERGe/eStmgYmMZemOBv1nJQ5EWrk8j1GrkyYwB+qZkvoH9hDqcZcTpP+HMJLQZjcIifkD
t8uwtbGNK+Ev6oIo42vgP/rsLx8olw7I03eR0w7Xf2Y9Gj5Fs8OZWxMpGhCRCR3OqqFfnqq2V3VX
yLeLn9IQB71AAXPrHkCBENKdzOJi+/1+yQg/Wsj0Y5RwDQ7R1zzZe9AoNhjlJ78hmdTy7anVjrkD
iWXwhMOHo9mb+v/gSXsH7wBGhIkQAECCB7KJrwq8z1EU+FTINjgJMZaUFdF2yQT0269zFAYJS3A6
bAXW7U4c6WdHE1jsxvYPsm4bCQxPlQbgXGl5RPD569zeulXBT550ef1EgyhudSUrj/hj6uPCthau
o3EzQpDT+fFDyTw+Pe3p9d3RmlJyIZ9ncH+OIVI9gIxAwM2g+hGVEgmUq07VTmkKHOj4GKreDDt4
O3q5kSbWVq7LovxlNkR3XS5mydof+jY1tuXwSzX7M9SzS/k20hZ6Dm82yThVdyH02/sTVQJYGdBE
v+eZbb62uYJMylgFdjqgkuPjp02xDk7CkoXuGSlz5ftuLdO+slC7c4TrNGK3gBaDxd7C4IlwLyBm
YotvNu+Qo7KN8R11v4Ryp6i2pH5z3/xzxwDO8gginggekCRXeeEBHxELhvHfHUfGps+QSk6XUIE2
PyQ4BMXeeu9EpMA6o9BMPhu3eGALhYkIRcYWMiztvDH+ClJ0F/TgzYBGJhf1XVqjAL2iPtUqbdMy
l8LnRPEOyal1e2Hqt47rNYPwL/qf3j2CLg9GJvDRhNij+RNwsK+5suJFSF22SZQZhnQfb3siAwVG
FezxmhVpw7rk71pPbQNvrkDA4cYb1y/C2To8KYFC+xVZMHn+R+Shx+qjKiVXRydSwaMurIA8775P
2UR9yIi8PlamfBGVK2an8ZlrgY1nV6y9ByREO/cn6nccXrgGZSbU85YB52cz48ZykPOoYHWrcIxr
8vXq9rIuHNaz7H8KOrOQfpn05MqUnz0EiCfKFRZ2v8WqB3x0cQ8TxjO2Si6yE9reGgGEkv8jCbgv
d/FlEa6iA0nO02VW0VjcTDRQn6ZfuGvJ1bWXzlCF4AA3sepXXj7UXLh68fRNL4vlI2jEZJmJQRsX
+aT5B+sJP8UutORBg6JtE4wwvWnYSYSmf7rZ+/ljQVZGe2bf3pyOqnDAOSbNNA08Ms8Cw0jyFtPs
/PCWFYEHWFs3X5O6AtqT1FIqwyDkomPOlVaFS3Vr3OtzwfHa7l5Iw18otbs5UXStFEJrCOeT9MQD
SUUggJcRbONFLamoOD0O5GXKSjIBSrCk8DKhsIAoadhiSCVbpNul6GOyqFsQHZy1Ebf/11XFohli
wZvvy4RMmkNqsICnP9SgRPdWxBNmYew5GOF3R6CtHQFjDmqy2GIGaq8DCkAzPi1dFzAIDQL4wuu0
dHFuzjroaxyWPF5xPDnpqvX8/5Ty/6XFxBpQoKtjT4VJ5kaEVUq7sqxe8OBfBKqW1fr2uLf6z/gk
9uInRBfokqMpXFNvzhLGfVTTTSmU821jAxVleluDHIm1tC/mcaBrlYRFgi0YoAttSeA5rx5HL/Lc
7Rrsq9UfQoGtr9krxgkOxSWL1nZrv5jeQrm2xMVn6sG1Zbjyfua5Dlc6Eqa3tf5D3sdCjWFi4gq3
RpAMTqP4QI8E2Zq6mUwj+vdORyCl7VzYet4V2W9T+PFHP6ULbso/Vph7/H6siKNldw93qfurygQL
g4nbhwGt0rqxjcDvAu14wI+57EHOrv+Y/s2DTjXkPPp+d5DxjRmI9vF6DgueCvy2lMIa2M/T6PcS
C/5LfrLHumAYVlJ5B3VMgGWLgXYJe3FFIRqoLSGLHbw0DT4ZKAs9jqSBWFBO0hYBCOG2/UFnfxZY
pQnVZ7bMVmG5sSC05XTFCj/lanG1RrymB7hnjflwEkuAjepBfgoluGTPvZpu2C96r0frxM292Z8v
UTsgYq1LBT0Y+ZOHjsrcOVJtTczhHBWQssgTuxPrQ5z2dX9v322yS5W3Bx/xIiAKT5zmIeED51d8
+mIeuaU+YqhM4C3Zrk1ecD9NKvIeeibD4txmlJ40NdEObLjIt1YqeipEF7rfwuYQIhBA35qTVbV4
VHiYoYAyvQ9BluLHZyp8NQjZqbv3pD+eVSoZwoSR34aTO+6++Og9d8PP12eWLRpI9QTlB+kVxhUR
0cBT4RjwUcqrMmOpfwXppr9C1L0Z66JDGC7VgOzFBTaA29SoE/9OdaNE97ITRSpMGFligVO4eh86
8/c2OScUAEgeeHzDo94z0K2Q67Jtv3p5xOuHARnOBB/Jr77WtMvgXnONwXLt6xjdBfeqJGbz1k8w
TNZJ5U1TY6VOrl5BQsPqaB9dNDubcG0+ovFbBTSLL6VUMB3slIBp/ZnoYaRwlCGZlsNckTMymq6m
s213uN4rvxR9latJJRkJzWlOCAPbjoUbRRXjujiROu27UioEPFWRP1XnDr8IzWxWtH2TXx+bDILD
NN6+ZLImUCN1/+8/TuLl2WMAvsTJDYYag3WJFlUT2BdMUu+Q8kUq24IPQG5yk/vSv73r4SyunCLl
JDtMeR9d+hb5633kCoU7AUTcgbHa4E9ez5wc2K3QYAnzup9qLp0P+fu3dkutvLasWVfdzemm6SRE
9NlDZZFV6iD9hc5Am0eUDqXvREBrzUhoCJo0GC2sDulAHkMXaVkfChnrD/FBDBswceX+blYijTbs
qFCX8loXkN1SLVPsEO+8F7ghpjzFPM+VTPi8qeYz4O5ahigdExzUJKw5Ri4VB79KMNTA+ss/4TOe
MWoJBbqfGNmaaOsijEU6ueStbzs+cvikUOVm4VZJybMaKd73EzZ5p/FwbA86cfqBQLwPm/5fRfES
UK7qDGV2T4oxDFx4YghmCsZPeIZc/nbdnIjZrJ3stW9th6aPdteWK204X+L5v3w4tWwu/C2JymP/
DQUfYZmsR+n+aASscJbFAthQRWLUZy08Ffiu6i4XqLL1yXASA9YRSZGoMuUcWOeDy+ryI1XYVf9O
q/gDpz8B/5vTxZ4QxNZPFlhYqzcgTInwB/yROcldKRCg70Usp3E0b5VKeNEDvN4O7tyiUtWiwLl5
8zLxOnNfqGVfJU4sAiErMC5HVZ6jQjgVqxs0Qz+jTk9SGYn1NFeDxagjSeTzLQjtguxEVx7+eRdM
4JjTLsCmkAZl6/BfmTF4mTa/ou185JU9jV7j6sV2M79m8X1FrZxAMc8vgitZx3j9/wDYdjvTRCzH
sBjvGwTLPyp8/p1ZkLdIdyJ7y8tiGT84b9KvBw/AvafUkB9yuOCF1KhkHJh2tqgnUc84x1LVEmD3
eYJDshkMUy33T0KyZFaLy790DQ1RsuU8pZ23IyLcScsCH4RUM28IJgme+0jO99xvplq4JvUPhtmE
K4Zx7TvY6PUrkk3MxFDcMVN0rUGmZ1g/yintGeKkINkNaqux8OBqQWSWPFMz/xeadt09+J7Zb1WT
TyjVbUFSCZSYLqYhJTQaFXc9L33EJliLUGT4+R6gfxEwCM0Zd+JrX17eNnWDNEW699vA82V8Mp4V
HDXwFdpZav5cAvEM0xcHTcCUor/OBUXLkXBf3tfOPAH0fBskjKIy0NGfi494ugvlhc7EtXe61Key
JmzychLdIyQWR4wiwJMqEnqbWtJB5ELpqjYMcSHfHr8Yxve7zzBjfnulg01KTeh/GhN5iDuS4Nfv
H2d+2MHzzY1d8Chu3ZEvFCdFer+g2s3FcO3rfQD9EGXWeRn/d4Sr5/nNlLBI1HbMe3/AZpZC3SvQ
29qb05R+W+xlop53jVYsPKDrwi1n5xkQ6TBivk/RlVU5Kb1SnrlH5QgMl5ekeuDUqFTWARDWKnsQ
vJz5FMIerEYwOpC1HgEYsAC6N54G+d+BERcfr1fgthtk2FbNW08ggBejKYUqk0bucQWH6SHSqaUK
SOGvas9Xj8nC7RGvbGPep3obRJkAzwDtpqoFXv3/pVZ8ozTPNi0hsotuQmC7leznzEwMO8iRKEJ9
aeAtUGqDRFUujTwmFuTl4N5x1dDb4LHI+X78Sc1v5vsixSoAwJbCQAUD/Q5iRWn+PDIFOl3b0LvW
zgBpNneTuX1iXRZOOHGhbxpwSHCSrAT4RSBAQ9gYmKZrvSpikRQupeJNxrIzdl+XlDygFdtW3erk
/J62FIaQL+5KcMtoDEDQQ42jl9ylmwjASOT92PNVRk+YznLb3GoHjEK7t0wRYorzCi3XNr/midFA
iJNRmxv30+YhnCgfJu9J4T+7Geuw7fiJS689IR1XD5IJMXkW2zZCqEEgszLGqoe1GN+20CM+a44Y
ARXEhn2oh1VqfMX9K3wzhB45aliItnsmWpPKhfnYemODb8gENlqG9vTROEPortO5njy5om4MX+MC
/kDB6Ayo4YLvqMegOfLdhIPvePPy+XweVAWK9ISyp6qbvzyGOcF4jPlDpjF3dJBgoHAYXdFig/JV
V4Zj865tXr1J54BeCWIM+J8ZXAGv8Yb2zUPlqnGicmJZsvKk92GkjOzMn76N+p7jtl+jHa5EpIlS
lEMv+2ATDeRs88+PyU0yzzVZKIr+NMIkbnxJvu/pcoyCVrcgS/qGaq0AHgek8na27q/Nko/MAOk5
MDC4kQNh29jcAJX1lvnemtgUDIdM7++nOp1hHMwNSvNc4eYfmGYmpaG89q9iq98G+f884q74MzWM
G2xhrlecF9WkvEIyr2Uhk/PaWz1Pqh/mVRvR07NNi910VeRIM02ufKR1YUwdUm+zjzzSr9Pjrdql
5laPZ8c6di62CAimju01587tDg5HtySqUka2JbmrNScOVWp7t176NYIsfLGJmZayLLjMr2L//166
BKADe9Ytw4YFANFOl6hJOLobNpXZXfgFUbepQINqrRsLX/XTy5sea7pcfLFXGVDMps/TY3YvQh0M
fi23E5/Cfb+x0tJM8qcrNEnNu9kkmNvJTf9eM8Nx2fj7SwH7nDUUI+xHDqECMvLlamxy5JYGXXY2
LwbJQPG27HXj4QFpovIgjLDbAt73LduKP+8Ft8ASuqcb+b5W169GD+5eei824a0G8ZCnMFauZWgv
u0jUMP9HOGnJMeiCEZmaD6oLWCJSTkJL4GTSs48OqK1LP12IO5OLRjenq73EOh2QXiUoIJRyyhUw
2RVjiRihGoK0RVUJ8IhSMwBmPRxQCtUy+pVFH094cpJ3YqPxRfyop2Awp62ccVhaEFyFf29Es50s
xZOl5Y5SV21xXf/J7f/hXCxxLwOTT7v29hiTxwT9q5u/NLBAzVZ/4s/wXsA2aXQ0MZyRCb4iKO6S
lY4VF5pfSBLhsoy3F0Ef5tlmzohdDEpYnFsNxssh+qOXw3sSK/Msz7Yv8gFKHH9RCo+bqzIvEWc+
hbrpraaKOzuy/a/KG6mP0IiW6pZEPA56v9mS0fseKjY6c3zlC7Nt0En1B0gjsG/QtqMRLvjl+u7Q
+cS1lBNsnGCATDzzQzGYzFsfMH970R4EYZ3NYPqLwpJWc68/RT8X/MSMrXzBTJyYrNz0XSiOpIJ9
0YKL8zwZHW0eJhx+lAELsJYbYDJog/GWrP6vdl6WlStewQ67RfkBOTxk/xsqrOZhIfxygSdwIku6
gUcag3sQXMHdKPURleCbmrIk4TetjLRU0QmRJ7txeJh9oek7LoOzx7CLvv5hSvxd41L5k7KFElsg
r9VGyW9hm8jyCaxd4mFDPV4zqoQmo8AMERp2scDaMreQm+xv8dRclvtQD64kg756bdJ0kUWuv6PG
SNWMdd9GuR8Tk1t1QK//jXiCIU9w8thcWyfeTDVANhIKdlgGZSGctqJxJkLDOS/MyQ43mOkTmHWf
fwjQlBDP3iZMxvXwCnBiltqzjymeP41dp2gI51PAvtGr6N3An3q/+ne0LwLwuNEh1WO/ZHOOQwFW
X/NHGBNkfNxPYcG047zjETdsO5sTrELmSlr/ySxgDHR9a0Meau7FgFI/1kaKkFbFwAu0xRqb//Im
tVc3TW4HCShtY4sv9BYhBCUkWXvl6pCFFzZ1S1Ez/eiGui1AUzX+QEaW5buhBqYNO9nc/0VPxkua
WRaSZKUB0jg/f+6a+OMroD/qpwM7otxNShVDt4aJ94qGPFwl4B9b31PkzKd3puTxTu/r6TbYYHkX
ZyS5LssTWURqZKMOPk8Ou9qQhymqPmfRlzriiGich6Nd8NpiEQJMiCjxGmV2v6fdG/r7s1jt4ssW
EgkAZ0iDR+J4HG6YByuid/SKs6pEu+Etymz6EUGfJuku/Q81awpiUKwuVlKOWCQ/tONR949yL58a
0J1C3PQ8zEHKLHhTslNnxZyBm4C2fCkOv9ICZN7o6BpNMxbnWIHGOa366EWcoubL15VDCSWO+9WL
6uyQNckZCatYpN3ND7rXmOQdPndO8D3zZHLisjvTZwnsr3Q0s/wWDO0BDbmFf+KqjXbxp5X81ezY
7sRFd3mehcHO3VZVzs62qgsxZ55D0LNIJ0MZWmJBwIMb/foErtwMsn0SUi9/8B92Oueh9mhl6qVa
X+D9viL8h9lgdmEZvU49oECufmIaoDWWjYb16K4+IQIFKwsIP/avIbpvr482/Soj+Ch4RYeanRBv
2wLJfc58ixLVmD+GB8LZ1evGvwGKbuiLQ/kTL49P0z19HJ5+CALPdPHpoZqdZy8D9w1NxVCB5g0x
u4wwYe4IturKFG3KYd7xUYIgd9/Bu1IOHW5jzH24MHG2pQMAX6ZP42znsWapfM5x3qz8G3vuIzyK
LGuLPTrc65GHJRyAPP23GQ3ofweE0INcZ0DhXLb3mXNDcpipLreCqhTXRvziPiLcCLD8Z+Uahk5M
UtaovvPNoNA12AE0R+khl1aREGAu44X5p5wq9zQN6AFkG5TlA3rlmsZQqPHtLXnpU4YpuTOoJzo5
FIlE8U+hkKaRGbOpMT764hh1VBjdNy0p83rAP1eOzSv0hg3dFmRKlzUEvLSRuRaosXP+eEupS4cC
B6NawaeVIlMZnmThb3iQl6iDF15pTmZ7xZRF7Fsxrp76z4swuxRjRzekgDiUHBx6HEWEUNkatTDn
uGr8tRrx4cMbxUjqbAUl4RSB9GGvEP2hT292kVnc0HbFbYc5LWMdpJK7ZblCJNOSEuWEqw04DXij
kc2vNaAA5vfsotjN5tw5iXkcC9Gx+SI8N7gD6TonvXG2pXljRGixjIcNPhDgyhCUNSwE6o1puAXC
KErIx8GFmBWo6pIsl21hOQ+O0KXpxvsU3TIxLXIUyu9cph15oyvhHsBYjww+Afzge1qMhdi2uRAw
2hKLEgcjnen+0KTdXmGAhOQSqMl3m4XEvFShSHgOu0LGZLGPTOhZoengL+rNna/t/XAPpnYhTR7U
5kC3jh3GRmwWtdiKUu+BVy+E6v4AARMPu48uSIyZiWBOVjJl5EWieZcerr931hauiCdzET13hjD3
8AtiXomy+ugBA6y3DlGUlqkoN9BY/CGixiQogOCjvZts0h/dnrlpmT8Mv3S5gCp7PqCJ4aNy3EQ4
02KJObwCe9k+9JgLuIVPmTXQWWp5U1+vtRBWatLwfhylXEvPx8hw/nZ54ETVaylUQRZi09GGljA6
DFtuY65IctKw98d24U7WTbHYTLUKZCpnhv1l3LlfifevWNvCCBtVWxLQy79cEX1b7GGKKygOnofR
5iAQaQQ6USwWfmJAIw/5w+uusqpfEBd3Tp7W/3yjRhCPEBism84BtCsTCljKRE6MDh7I9oLNl9Za
G0DmqDcSgF9rZsX1oVoW7jI7DHsjIHPbZW7jHYQPGzovN3cL1YAU7E2r17m+ybk+G5Ti3TxiWfsM
S+GMiae7XYf+vrVnOT0rDQu/AfNPkv2T09O+yDa88hUQJHktvw5DDCLulMRsf3aruBbyVc50X6IS
GRThcefYXbycM3v+PgIwtgZSi68GOqLNdn5XkJ9NQ2LiBM/DHLllhYVBVI2ZNwxAxsUgNUC0ysFY
WiM+S+DJHvLlZocbq0RX04ZRbHY69HOQHEC0xT+yx/neRGX60sMIHEPqAjuIp/uHPL1C1VLCwsfz
33lnm4c80V/D8zPvl/fw1UJioUVSbBZiqQkfDvnKPPLBTapGApVU3J5WIn8Rqsc5bSl2VTTagvWa
AJUHbY34+JwAVOvAQkqQzf/om8zfDcfjyrfoQTrK7jjOZmMOl6LCZ0K+Ap3UJd8XgxsaLv+T0iPe
N1p7J5XEnQgQt5IIlf395CEUbs57e6AKxR6PqKqt4ToIkb9tqBJxfU2ap+k1jdGueTTbcb1tHFQZ
G8HqTIFi08OiMFB7LvH4Dt7YGrnVRMiNitSSndq0rhmmhw93dxWnenUE1gBR+W/iAblzB2bMhzkL
dCgbrxWyBv+NNjQItpyKGJXOxisEJi+TfrzCLJEyoNp11OJbBxjTpVov1uVwJ4m3pnunT8LZsN8a
Rm4TbbkTnhhfw1SMulDBP8SX3RlPx4j6u0yTGyrSkXhGcSWaAWtsmLzYq4IMddxyvhbvgG/d3GW1
WnEDVOVbz8DbCB2y6KpJkfR4RuBiiFdvoD087YnGb9ThB+yHuUGdn/VDN9LSDI30rAv0lWrswWff
oH11QwQrUnK1upW0If0AXpo4RckqlD4QnuNtCMl+/FTTN2dCSHxXI2pgsHCWNGqRP+ppItRXHI21
L1GNHZEbeYeLYHqmwcc+QxlmVK+34R3X1BU160gdKrgayIcStvNsp04eKxsYHWJoGbdE9pds5ovp
QB0kCGde3c6IZah78hoFNUeQGkxyR79e5vYwCUjOrTSJNNZvsRG5pHw4P8D/1YRs+K6KLQnJXgJa
k3reS9QOXwOmisz6KV3O0Vq7Nc6wwLVPnP0fYFE5IDht/InvtyVwhTMSVDtSmgvy+hAgNhQDU9mn
VlTS1i5kyWHEm+6phHosQGuD0F5I8EVFHlhl/+7/aMS2LF+qpsYVLbp2J9DT25MWWjCjRu4jXw0Q
BcJ7nS7Ezpc1tSXFc9GTJcgZOjghXKL+REA0KArPSOuAcMWNy0obd4E0KbyktMFF78Pxh4cjOCka
7EnGQ23ddeDRqxidFsezcZ4Ty5rBtlho7lz5zkYp6lwN61IkmGyKTMuDEQLDuRv4P0HGqMU+DUI9
Ib0xxFc9ubJLmC74bfzjHUUtAS7ubRE/RbpPLSQgHxvXQ21MNeVH0UgidNPUAbVbpTMa9tMutEJS
lPX60xpceuKmhb///A5omkNrtvwi+n4uu6ZE9PPbcJF9LYoNQPz3SWLahYvT7g1J5W77aHOidlu8
xFOQDVTeH01tGoH8DTqeB+sen+Xl2Y7nvsXJYt70yK8eFmDz/4fviSI4uUBUgnfKE6sITSGFEpyR
aFMk8YotT+EWUa9hJp7iDCbm7TC7itRsJ2c0HF5AWiOyatWKZshSZ/8jIuquCt924VzBdZIk7Epf
zHNaXTwqFekvgYt1jVXrjQy4HF8jkn+ZF/8N+mA8zg9W2w8EzSdA8dk+R0UtpmhElUmlpXvg8s+q
s0r6CFZcYw13nNa5uGKW0qvS6f3VZxKlEC6m7kqo0tALUAOfElUemJY8eQvf17BOyikNwjifIhnC
2jndrRK3wrUu70UU/IslOx1T+0jSSJ9kW+rPHYFqNZtfQlaWHGIssJ4drNBKaj/ypbnZpW9oOcNq
OKaKicN2YFPs4s6R5s5q85FVrMvwZPWWh2R+Uxvis//xRT8Phfrr9xiTpFLZ+BmmTjIsO2zY5fR4
ROvVUUrs0X88upGFPFh+53Hf6ufJaw2tqQfl07BAOTCSSHhNy68jNXIgfHyHVY4E9RbMttL2R28U
dD5TabgZMLqO/UxSUIIYJFsRrJlDs3DytxyOM2jtOCaUmuXpYvnkz1LYy0bnGAQOCIYIgwPD9oLB
RqKojeWL+eFvkvNVhvvbSJ6+BfZ0PXBZsm/LkGBnxEU8S9syFuxnfxgQPQty1Pf6T60G2+BzS9uU
XM36GfNY24vBE8r9jBjRcfntAwgjBvIVd2jQdF+PU89KxjzhhDDg65P8TOcLFE+DsAwmViLx6qzR
//Zcjp6iWA6aIRcv7I6xMiOIvuCud7SqthXx2zc7O3wwksor7WQkrmWf53F5MFjMA8KWIeAz3lYl
sj6v+wjlYZ6Pz6zVXtE2i8t09cNqT25+Aj8pQb6t/EMpxAszq56zJ+x0g3jrXZ7qRQeFs0Ws9cpd
ZZ0jzDRGDS/Nl4NnOqu4YFay8tsZnDQ/qFvpo2sefn15RYhU5rMKVt0NJL7GKc+TPIgwnSH/WIFY
87sKGd/nndnqXXE52zhaq6yiHDqSQ6a5bEPOCoYRc8n69pdEm+TkBWvDmTAkpTznLGHR0B8a70gB
5usvhIwgaBjj6UJAFazOWEwofHWA9rN4jgJetzJeaKoUBJ7S5Z65Tk/fb52NS+XDPMeUHGzQP0z6
z+BO9vZ/zHjKQdfeyMNpo7GRadGoBFLTNPbuJMIE5ZVcSHsczpCqBk+1EQvkdbihFmZye9vW57vq
Tvmm0G9W/3otJJuX8kTerIZxTjAz6e02+413vabvMRw1ndCeA9TSmtJbkm3xRFpZOs6BUeaefCNv
6bh30cB/RH7tT/c8r+/NdLC5gfQ0SFdxSOs/eSolDAxgBd/JXDH00OIKCQyVy9vzrMS20E57p3G1
Cl9/vP4QOhOxCvspLgCFym6y6gwx/koMeuf7glPHtFsRFgdiuL96GUw4zzreT7bDUySO/E4wE+IP
2ePSXxtWK808lFD6QMPZdNRHdd9N388SGuGitLhKlV4i+WYxBrGc8muR/EtNfM4XQrU1fLqAT9I1
+0bMXWkGBflShX/dvQiwlX2twxEeP/IMphNtMtKPh0tnj5zdGGgf9dZHBsJz8HnBKfEwC36uCilN
jDd/t/4PkjKjRNm+R/9RyXzG0zRwe0+SQ97l5X29DUSKHoV+6eUWgkU260sMj3/6Qd52zhz/9yDk
lL4PsKGJiRYcJUY8O/4pBcl2gn77RPKygyNtz8xvQdZ1t8CbZYwyeX85Bx5fMxFbXO3orPw14jVV
meXmj6c/xjJ4+tAZ7LZYJ1MwwKRxfD9Y8nXZuDe2PQ/U6UnDOob1RVvQqx4JlGgb7OfjKVxaO63q
103jSgu5w/C6HIXcAqFoKCEksb5TRihjFlig6jLQoHnOtSCKFLMCY4qjJ23HMKhhB6xOzTdy+cvF
LmPmiUF4aqO7SDjyoXR9lpoRezn2HVIGAfrLdZ5QvWdlRtoAxWSEL3J1qms7oNWNAy/kkvXj7CQw
UIXV68LPB3jC2Rf+aRT9NMU9NwnfhjaW/aobdu6ssZfrmw1Vc8f1BimxRAgvEEGjP148jInXrq1P
MXwSlx2hXaxI7GbGciwYlzEw+hwlIC3xdOzMKZMPFkMMTPfRz+3by5xt3rRqCMnjyeKxAIeQObqb
fIVThInqhv3pOp9MFZkFpxYMT/RRq1nX8JmUTLHvZ5/HBBzzXj2bxgZlWVkMb2C75+VJjZRUstkm
nzBsT3LppBYRt4y+ONDzqG1G8kYv3dhv8sepOIvs2/S7E3FukFXgFfadv5scqR4pxBCqWRX5E1eC
9Uw0rowQ7urjTAioiTpy73+Q8tWCTwq1kFjfapR3les8w7GmM+aY0u9Ojdj3DmSI4b/sFFQuE16K
/K1LuDIJxs1P2uD0jATnpZ4N9JhKFXLbEtQst6V6CLKHWqxpdnCDI4EOOBMtOcI5Uj4Y59etz3lk
e/hw/g5tdVH2V6trikPVlP7MeBItNZpvvaqabE6mRUcVvNMO/fIT0FXHtYrTWzdtxj/aYvXYJFEy
28t98BySUu5mWmsetryuyJjwi+zWCyvReonl4PZ+wWdqgG1qqeGdt/uvc0wNyXq7zuOUu747SbhK
qL2nsqTnTVspZE2HfegUJhVurUqc7yUdMzERHiKzLmMhcSwO/hM1910f90E4RiTLXFgF6/qsL/vf
Hn1kJ73FqO9mfeh2xVOjhMQ3mWn9Q6v5yTMzo/jzUJQQh72MPlwcXM7wQF68z3e/7P8rcBqe39aD
v1TFEmRUbX5ADPO3VBFTRCnPVZqJwHtPCCNYV/lWGjLjlbpT8kpiTbGR16LKDAfWgPvQzCdGntJ1
wv4belIdGvA4RgWWFekNwpSlfIK+GpMkpnGMV3ShtTj5ilJ0hS+1Jfxn+IGDStBzu2c0/beX2gnt
p3eDnuE0Lsd3GzUwMX1qf2g1xCBmJpwwUojIeupU65n5gnDMDDJQhWDBDoZxZnPXdF5oUlsWUL9M
GHbolxw9y3CQlGuOYYhpwxE3ZEZ63xQFqkdSYpQzd0IL3cJ+5cad49IDvrtNXI4JiM32c6sH6HeG
381/dHAcwWtO4fYgSr7KNX1B6eWMy0l847cAokrTFFbVllwUpKlxZVtjnqiQkrXSGdmlbi3dp+bD
fVxfQd0/fZEK/mxvCfO587oIsFk3I1nmcMW3YbtTU59S4gcp2E6QndwNMwR5od7x6UsH7lffv7kM
syVB7bj6p2XDf+VZ4iUcYZc2ZtId3xZ55OIRVv+a+WgPBwkbiTXfgs3Jp9yd8vsm1ymAST3Q4gU2
P9J7amIy2gFlFkj1C7istYsnbRIvCvP7i7pn5/NH2KXRw2bL0bCFOOhl9n/VIdWcToZP1AC4TRzD
0UD0EBIw4hz1aDsXqR2qb1Rug+lJ2xbaKtHe8sClF9iomD5OtI5toiiJFSicw6cNloRXOnuNlOnw
jOUHxHsr4KTG8ou8Nn24LTO9zQeDuGLXfNEZW7cwQdl/8kfDjt7glq2uTxRN0lzbasgWkFbLpISU
ERHzddiTWLqz2LRPcMlEJc0u6mUBCBqBxirKBlvL1k/PZZl7s87lmUC7CY/s0pEzwZyVeKIdBAaq
8wayKcoNylUOKBV6FjgCmxU4PkPVVB69t+IX/qw6QMp/7CqbkvlGKCCzLyL4D/VDXlFzbpLKS1BS
W3PM5qvtHc2KUkSjA8H17Ex4WxpQV/8ss1HRDSFc8JTVo8eTvg+QFPhHfo8CqQ2gtXOuwiMtdbtn
sHlmP7cZ4UMdbDWQg2/YEchdzMbWRrskCM/PIoF7Sj98S8SgTKKwwiCxRnLfOJbXYEC1UDN5T1Iy
desJ+Nb0XmD3pqWWFhkskFO7TahJOgvMGbRkSr3a45gGupOVEWSOwAcjJsqhsMFcyeT045gfKOqn
nhKXrzUYthDeXcH/vm0/PCGtdRxmS+lPPQpebP4cEQyDpSSZqm6jybkBgJoIC8x9WgOzV1dndYLM
vRAQNiAmn4PjVdlA15xVtL4xn627BTOf0pMs+DLrUI3YA80u6dPCiyaC1YcAqUCkCZQxmagcYwqt
vUEw+Qr6YFzO34Hqfhw29qQqJrbZmj2QvPdeYEdU3dVYT/qgpGJ1trwSWqealFt9rKxyb0HKJg03
Wq1zpMksi2h3ZWF8EMvLyNKXip6dpJyyWNzdF4hHtRUgI22bojLXKqb76nYWsnEmamUlNRwdruD4
X4TjstAorOLfY5pMbM83dFH+fQmXkDCwYgTdPNQw/qKr/2CYh4fJ809rcGQ7v34E+PD2AG41VZHj
f/saNG+SiuG/2e3USCQcnHhHGWcK1m2pIjKfB+FBfeyQ7GnW0gC730nHp4hSf6ktsCGjnbjCL4zV
oaF/kiYLPlNVFoNE7+8v5EURAN6Z/8AUU+9LlAiHmub1GVuD/Ru806/F9wOHcS1yflGpNqV/tHGg
iNja4FS2dKvtOtTCulNdaWNjelIq+in4fpTqYd5ynlCwdpSKyZWr1LV5hfAYPnX4N4/WV2uUTkrk
LyDSpkfCP4fnlUKGSyVl9Qx/II+PrupUufrcyoKrSL1lp7T80oKhJa2IjIlgtE4pnW0WT0UrkoNW
GzT68EObqjDjEmTOyKE5y7X3UVC4vNvazTLiWXNXsl/D2kn/uihP2Try2OmiqIZJ7e30IQCopK03
IzOlpTFb3N0NRSQ3gsZ/OoddNlsS8FlrPurYSjBwWe0NJPKAHJzFRCNVn5KbFA2fNOcr3gbPRRQw
kemISBpKe3dJbFcs5faOfSn1D90TpzcWic7Mqq7SZ+AaXp0Yc+34NhqSHegDo3dca8dOmbSnj975
NEVdrxDyfFdu9iNPFS4aOI9XJbJk0y/8zn0g3UrZK8eP37hITWD+kKG3yhUfBfYVOJSyjGs60Zjf
2QHMU3Nwz1D1AfV1AZUTFO48NcRuzfCeW8r3Tr9ijxL5R5VmQImrHr2dsQMt2mJkZ/Dzb8vin1+x
1rF+fOm6cm9avsV3+bcpzySspgknXthEgH3gm4UuWwuHAscy748jq+pwPH2yiEJtU91q1QBrLc3G
WYxd8R9HsdzXHCA7LPp8KGLh7cSfAiIq9CRrpNKLJRbWtd7Dar33kmbM0qhbHEI/4m2V8hU40d3a
eRzhxQbBZbe+Nrx6JJIk8fIfsiJlOM1gqMPItIXTK/3b0gLH8tDnrTGoM/zku/5i0rhQmz8o+09f
tbotyyN1A4bNITdLbpde5EKFjksIcB2Wm4z85XVCwrkC5j5XdWDq0FdtVWh308OZDCUfAoBkgWZx
h2GM5zLsQP+o7wGHN7gKpwUzZEcRYASm6yRt5JvY9Mrc4ASGJkg4yIHlfj0yOg0CNtyRk3wf41Or
1CZMklorGSyrEpAsp0RVnQrp8yehn3LfaYyFB3lJholLX24a6T49x6jI8QqMLG1E6gg44rzISpzL
WXVMqVOiNT31zsm5UjLUzcNbd+z/aODf5sHJE7jXUlBfmzzDmzgfAHRaAV83ULaiX8MJUKTvpL/S
al57s8rrHP5MUpmqrH9Nh+UX4sJiTdVISD+WUpgnfRTUyRSA3dyFqn69T+kC3cQ30ilKqOhVQkQH
9fKHuw6SE6uHOMH/8n0PWVgkQ66JOIVJtR64J9fzbtWnw7CGqRXlNPhxewpUG4+znXy61lT71chF
YXidbGBcoHnLoeCdhYf39hvYIM+wpmoDsD0EnoWfjxwSuR9PqbtJHbQlyX2wNggSnTfxaVqP3MsI
rGmZxwiqXsban7Rc2joUwb6XbwgSMs7CKkDhI4IgGqvtbWuCT0SEA2izdmKLk8A9/xUOCSCXaUZx
hFaWsRbOTmWnaCw9uV+BdJW7mhSBZYUJwAfc1tDPiGR8gmm9Qrj5F0IMUbPKDz3U9qsLFyrgjBoO
FiJToCwhHmTOp1ric9SCNR7olfM35T4LHJ+/JSiGL2jjIcuPDoJ8UIWkpZqrY3BbZ850f1m8PIYE
wA4+7TxDOVSQYsRl/ZYidwOkGmBKMGxTv2fCeA3lPOWA41oMFbEcVB1bWiVloHdWFp9P6xe+AMPE
4b1iLgzo6mw3sHn/zu1f9tW0jNhhWYrxKoJv7MVP40jUN4D6DYVkwzPyQBsu2I7A/6F80IRdwwKC
FiaJKzT0V/jE7Ptj+r6Guhi3Es2HjE85cIhYiBWWx12d5Rmhq8eHXMKaCzHIUitIspWsVWFv8IQL
qesi/Z/DQv3yfVhXdGF655JirKbzlzioZRwZEXc5dI5JBddJqlBkfjRdSSJya5hpS6c4o1dfRmxh
ckaUpnl6WjXegx8GU+tee9hLRLxBYUoQD5p9/kLryCS4SzZB/x9Y9EbP2FAQJ8XrziFGZM/ReR8U
comKfVi425oKW8M9FPX815GhCyXXC0G/0eAME3X/s4YxnZFxMBoMfujJZ84eSVTaNXSOUyUxh9e4
O8YtuiKHPBmGL7omJlWRo6hKPv5CO6MixgkG/evPrFoz9cFXypgFR02N2YZEwGPknFqGzu0uYdtS
OVqjJ+06a/oeg16qVYRxzweqe4WT2cIf8VqqJ6cLEPns6bhwinFY7cQrm/pxlI1RUk1HWYnNPkLa
spLO0OR7BS02BVJm3b8Whj5aqlGcPFzyAy6eMbdu+E1HqmDnoFT8FIA90VZZV0rcQ1dRN2qr0mD9
qQQ45+XyRWDNNNYsIw7N27MpumMZ2O6yKAyXvQi/y5HIMhYPqo0EwOTR79K+9rFl6EqM+KpCased
Bqu4v1tfTDqDQSzTuqixSGsSncVW99g+Hpvy6GOEobfrvpPrnR/dNgUiU99O5lgxuiTPd5YQfMTX
DeJaXbw0SrTL5szgzPkQVuMGPPJulBBn9Dix04Qall38wXZNp9fRZP4riBOZTQFlGq2aVhxw1Xr8
VD20DJJzzmIPlWh8Kf/fMuJYWkAxj6PvgbLquBxAbbohsEHjViKaN1WA2DqZ5A6PKYzRfXftb/Sl
kvHrUf38FmlTHBBIE3StM5wAfGXfvLCiXfnsRhncTySLTM1YkVZhC8UFpGLLJQ9pqHrNGsiNphjw
crNi0Wvlk2hdSeXrZm9wwETEJbxIvpHxnhFeCoKidHoS3mZD6DTnO2LZEMRUpPTtXR4VmgA7X7Df
mJQgnRqG3y6pfT8W3hxNYX9IOBtQec32Vs7hv8ILwCjr9dJFmEKiFjXy7kPrCYJeSwdO5IJGPX+I
JXAnyYyZcOEx2vbyF7r6WNF1a0yrrRc2IH4BhxuNT8YGf7BEtxhi3k/dEKPgRB+WzzYu/ktZ7Hs+
jYH+aZ4OSj7KDOlYmhHPCk2mzRsGLU5nfTyIzJ2HKJOGYtthMugYiiqapiP6APnpirSQ/VbSfQJ7
IUHUxTtzerU7i0ww9s25VO5kCSQKbBqw4x5M66r59xST6WG75k1JA+5+SAOcdfwwCOcfuBbyVIlK
EBtO35SUE5xIQ27DqgGsB0eCkWm6tLd55corVQrD+r5z6eMCpt3NPRmuRvIcDsTknPQyLJgdzGXr
NxXp//xG6D3uzRnpJC7evyua6D7m6IxhacQzqB2vW5ZceACdg/xGPNSPeO0qVhgwA/0MnO+Bw3kn
0Ak3EJt3xr2eetmZ71rDe0T201oXU1EjUDtX0qjVhjokQi9b/HENAS+rGyt3GZ7WoQzXWMZl2Sos
KN/R2ZcuL9hogqi5BfXgPK6XSqiqsfmRaDmpxbwEnxbgJS+Jrjh1mZGqZSa/qhAv6gD03U8w8xIo
kGrxHuE81syf6WhCY/gMiQqlQggRfu0ECoT2YtxYxwmcGZKwAmNwnwxizY+QmQVDV8VPlsAqYrWZ
67SLUMJk7BpiZNqsXnbFJ9RuiivWHLH55e2wC1lNZRSv4PgRHGM+DWEOcc2dGWWCn9tE0PXYqe8D
wxOldc71MNnLQ+c8jbGDX/IKdlGslpaqOHIZGUjmZAJGR2UhfKAmOtn1ckLfPuN9G/55XwxwG0lo
/53PLUYk3umEPhZpVvGyQX59WYxSI1k/3zPyff9fxMCAwjpxHrH4JWykXgHl6J75yLRki6nJwvUs
Vlr5YdhIHeaiuqsazWGozsj8Am8G6pb4pfEXYnLQiEsC9nZTpRzhGFmpZO2Izw2MOxUekSISs/Bz
jUKIDwFkY79tPrVfae2MA2O0eBPU5Uaq3Vz6fHG9E50PrDxeRth12fxF//EbdP5cyfcgf74jlSzd
ryy9rnvVrDyCsozxO00c2m9O2qwmOPTwhbDSUAoWZQhLgYIY4e0HJ6JqHZsLq+xCTMuYxy3yYBFV
+EqVgytljHHQKizHXTvEAyWyRC+QjNyouki9/KoPoDQhFbGswK2CCMJ9G+A3HWL0xuo6CnyYOvTP
OHea7vW2NZ96sBIQdG2HUEO1Xk0zJxspBHkTMh/oeDjS9S776pSitIBIlQnF9K0fsDBCIJB0ORQk
1dM5rvJqil8QIHmlamsorc9E3ohEPx5a0YeW9Z5Ln/BefAIFz7p9jOgHA8T0MZVq1zJm+fz/DNDg
LpypNDJcSxeomQlvQLg9cA3LzV+YronYsWeipOhj79lA8pHp1x34zD1pM4I3cRwCzICbvpHi0fos
tDbuYqzjUtSH8DDgR8JUTmKYjqLIb5RYK1zoIw7EPivOX8/EZ3yPuvpb30b0kX+WbqqPtyP4GVWB
3+TysRnFSfeK8ETe6d4iWVjaFKOfIGsNhLPV5M/A8g8RmrCz4lDejoYBI+WQNfDZWxK0nSGKc/BF
rGqJW3s8NKH2Sf+/ASVZynIgJn5YKhzkJibofDpZaHvS9YUANczPqF0uliijwRGCqRpjnMBa11NL
hixqkAAelRh1wRITNFZgNvfOJgVgAJ/QRxrD6mKYQxlt8RO+aVxTMTPzeIg6tA4nlKcL5V5GjoVC
YyUQSkwob5rMxOuoBCZ35loHRPzw6MQAfTR/KCIT9UArBmoxo9m8ga36GChXcDkHOoiNfCt3QuoI
JsGzzOWNriNPSlAIxUn9u247i+pYiQ9lbwAQSND6MAZW71Bsv/8FHZJFgVqPG3FsWnTeGBuDG93R
RTcvH/dEIAH5nQe0NoUlNDi5t5QGjJvpQ9KlEO1xPhk3FUhBqRlf2QJ4sDP78QgGKDva5dW5+z2K
XjV/6Bs1tUe1PqKGmX1Ef2ObuLUVsnA3nJzQM1quhZR30cwYJfXomMLtIBP3Md+RO+gBwCruK8dx
XV0cxz8iyQ+pDgjTTzfjznNorAsPJ+A1P7W/CN2CO8VmCFKN+1lBCFPg4kB2jaaGPtFpX/l5iOfz
BgRJ1ELHU7YysjsLC6DOpLvxzR4G+dyUIgjdH0WHyMbErxGq8728qjDdyJpo/gabr40wnOM682fb
GMbPJQW4Sveao1+683Cm57PRYI1Y35WywKL48w6XaW3K2ubXbIGLHEIkxyvPRC3jTrrjSWFg2yV4
iZrdFbG6+urgBHBFmjroQBNs9gvGvWxADXnp/2OcFVIXhiRdtXogwmhCKPQiCV8DtxxfpgooDEEa
ySddPvcvHga8mY3Wkd2qDZ5ZmICy/bZJTEYXvecU9I1RQTWSuHCS2fxy6yFvZIoCVM8NijttIBDz
YvflJEU3vm/z6tVDINBSLufMErvGIRXJyBtXCxdZ8/v7bjjL6K2vz4zHqRhjYRcKdJc4p/cBLyyo
4jhgDu5GFTubYTI0LpVmfppz23WmtikVCGoFh5vH1aiO2ny8NvEaNutrJctVESGNbIMeh+YtHF+L
3mo9uJPQBaGwQJolM//evHAHyHtcjxhqjW5D9t3/K3WIzqZllJhjVD4/PMUX3QL3pe4/1UCCXsam
xGT47nryl6iOvbvQxbSrQPNqBySs+TWgOw16GCiCm9i6WCPhjsU1Hpu8Ci26YdtWyffWJrqBVrKE
qU6/JULs3J5sPjEyBofVolCYGbAEH3LrMGkfhv9Rdi/Z6DP5BkTYHKh6J3A//ithTkaojZlNJNzt
AMbrBDHQEbOLVdBv3/69/XopcN45Xt1ksMxF5iubzoevZ4hlNm7P8qHZwpNpKSDlcWvryEyruVrQ
IoMTFw9QtG0Qv25wt2UIblci3Z+OwOnzcejUjqhCoQ8LI818oi5ily3idbmBsaIn5ww+gPP5UAXr
oQkqlWvL0g7/Jssm8Fd6twGr6g/8lo26ABrb5z+CyOiuYXvw7Thsy0lCyfHsIfWnz+h1bswxMtIw
7mrnPSvRaXtbHRdDR/1dNASFQjp266vwdaaziOFV+6+6TCJT506vl1KoNdtb/vQve3KgY02loWXQ
ne31vacGPGsg759ni2eIQa3TeRgKCkyi1xOj0+QM2rCWzAQEocEqaR77MQRj6Zs6KTWfmAF4wl4X
SnQDdU70VHNKi4586Oz59NUK+WO0J/TnY56xvj/1JQYhg0mLNMPMgJHiW904BvNn9hNH4xjAMHLV
TJYQKj7rK9+ZgmEm/mYzXsvV1Arcr9JU//yvg0TD9tqiVNpGOl1oPHzCLvno892L/C/1mCWSNc3f
M3TQZ29I1yf24qtquSRk5gnl591Ci4ZQkMH/ndP/8rtFF62CGc/IL3OhtgIwlMaUULrXHuA7b7oG
mwhBhopCqZFjo9yGuqsR/gIPwM8a4XwOv2jq2IorYz35j+rna9b3+WDaR/stCuL6ixYZLL7zqwwP
jSlGM39Lh7/onoXldq76CyIpb/2BLgYjlDnItuBM2+uVoTc1aBf/s/fWQv4eIJmH0sxWjkAr6GIt
IANLm6Q485GTkcFsfM09+e3OMgtb+huFMG0P63kxrVgTwSbWKlof12jDk+a00WMT19kcCotJ0mix
6rZIWv8NcgInfg/1dr+b24vGH8WAgd5OKXjM1FPwKidza4Xse0VRfdrcGksS4sx7jd3aXRFb87u5
Kw9Ct9hzOTrEirqsHcRBfIj8c/XxCdV2nsPavxweF3WglUGxnKh2E2MaMMT+f7Rm52npcQcKDzK4
ffVjV/BounTZUMQ202nk2V4apOjX4nemKYfQk6+T7RCGl7KaNIucry9/NzfqyVhqrLTgZYAYn98g
1q6ozhvKspZlq5S3ebLTz+j06a9cumSN8mfu7j0dGRbp84Sod1Ne09RchO88BFAKlCDpi8QVejZS
h/K/yv+64in879ysvZrcG9rgxcHhnJ2cclR5rb8sdXRg9lgFbm6PHn+hZIQFpw9g9U+UmEy6uuWp
5gXgu0Ro39RyB/slYx/V2h0sCUlELPd+ZHH40D33lRNaZi5a4FEMyZ1/MjJZmgwU5ZtnHxBPRFTn
27Xi/PsE5iqRzrjNyd1hpaGvDir6AsAdgbjshCxO5yT72yWk0fibOAiKWWQZ7X1yHkzM3dvjmN1Z
FZKkCohSbYb39j77am6Yfi4DQbOp3+Bw/AYvVEUI2gCpV/nAf7CXS3qGO5FCimTjYiErPmzz2z/v
SAnYaPXWC/XGGFI8YdgeYPEHU7FFWgkayrT7K38sOv8iznMCO/bgsdiYPJXtI8+5GzwAv2iMaNRf
fKEc7MJYl0ewcN1k/G2bnZDuGtUBwk4yJZ0rBa7nB6jgc1k+PIlhwyKN3Sn/SVLhp/SNO//p4cc3
KsOvcUAgaJskiEYvLndoTXId2jIvDPWSzCv9cxu6w1AtfdyTHoDzMlQhdjUBmCtoOaRxoAAL4jRe
tNh6w9j8f++968BNLxWXxVmmIBugkT7d2urcFvCKpe2xmy/4uXRADfiMUor+00IAFkXgYaDAcjL9
qIDQv0z9qVWn55cIWcpZHWH5M3jbY8ri1OZybA1xIKJLSzwjJBEuVW02WcI38pCArHgVPdfSDZo2
k300ATOl4XEDduXZ1of7rZXlwx1YsYqEKJBwJQdni0WulnQp/V9p6l7zR6pcdVqLT35MX9ao151p
gHn+UXAohODhCg0lhgXB/6PmJEokJhP9LJe/lsbCP48cftWyCEtDQh1dsJKJK5/4RSfa+n1N+FJe
pI4rosPpg/BX5iKSvANAOo1Pct17xqfniEHPdibDgl6VemzpGTgkVkTQTdcS+dTrVU8Als5RUqEe
JLMo6rWLX2lYaRePwneXTmBHpUe0RrjkbNakg4k4N2M62HzQAcu0AqJ6jUzTwGLtUjoEJz6G6WFp
ntixDZEYzQVqDFVzc+uFt2muQqaktB6KLMZkR9Ndr6pJ4jVOoZavgzUAsUNQ/USGfuWWGyvgDyU9
Y3vbseYvITlfZrbmYUcZ2MVMBjuqKTGiuDnRQd4DXhElXpFdh9lni8F9YU/TPJQExRFO8bGeCFK9
cf4af81FwR8/3Gfd4gQx4vDG/1xd6Q0j3cBAOSp4j+Jey85p+JSJvkmIta9zqZa4jVzMHe59H73m
3D4CfQ9FOLBh1/yPFhezLf3FR0Q/jcA3gChgjJbctlpJj8xV5GnkrOYkWeWCaZi43cwUQLaisLCm
x31B/Txsk+DIpdI+NCC9wGA+K3vE2DEgZg9WgZAo4fBNUdVDShYCHC2OGIk8KAgZFwrm+U/U/QyJ
/qqLCEErZv0vbWPQQG72YZq7BSpdVlj07jOovYtRvZl3VDXaP2x9MKuPdv8Z7/IgOUsVXV9dBWa4
ckgZBB7Jp9vYCJBfYCSN0VAxg8LgVoilPctZ49X6kcvbxA+VrJJUgnbNCEtznZUQBWG6Bt324erN
DH9twKXIICHg+xMk0x1m75fpb/aVzfHg41ObMD5mm98aXOGPRDtA5nNeSM3ICo+5jIDDSMbbYAIu
vntANthMDw1kGURLTRuV7kjGRfVqN9A8Hlx/zmy1YpBbhlLDtVq2xwXhM4o73GBNOovItjOY5S4j
EHv4toB3/zNwKxcp4yVTopjPSAg7PqxcDP5cGUBDLSdNHsktONo6Ctk1aE+u4xhhIL0rnxv1gKZ4
PY0jbifa4TemQvFaznXLJXDRjg0wYv/HzMSZYgDY6+LeZBeQTtsKjCtM1fW03UZUl5HQqDv9suDK
1miJpM4UEjUr9th60Phv/ARQwbwZumMt3xXG8vawHQge+gN08Lv8oeYIrl4cRU7CNx6sv3SkVDLg
3fME2LVhCs5vOlIXH7vzQi/klwezpGQ6QFnIT51Z076RT1VANFP3RKOeD04RBjp9Z6A2rOUNLD/Z
JPgGSinEohry/AScMkbiAwQlCRYqpQwBscUjGZewFLwD/wr66Fhg4JUby2WazI6kNajj7SO3EtkZ
AhK9OxO59G4MG9g00/RVAyPVuEeNoZicZLW94vIHrt82NbLXz+zT/q1KzUy1ELK7wbzrUCkiGDYB
znGRVVxylM1IbXbjcQzGqGIQrwJ9DctWluKpzSP1FrXMDM2TnENyoRivVgPOcHWMW3zK+Yruo9/B
OSG71L3QZ49lu4nUHAtcAFh2g2sVH2zb1FPWEfJ3OO22QjdTCYmD3JjuYYTOGtFq4FWlPU9For7f
j4Z5QRAr+z+E07h/BrLZzkppBNdRVDrLWAieZce8q5s8ax/ZYzTojjlY6ABl8MAXXIrsoZc2TNKd
xJrClZ7uKDv4oE4z20lXkql0+FvIaRxe9s2Ksoe4jznO2rXU6hUgzbg5jkJqWccKWiS/9kSpI5zN
Z3WA0k+QRYTx0ZiXqZjGU5zc9QA2nNkscbbAKKgwx7kmRqhIO9I1hDGeRW9v5eCX5htURgvoQEKb
ZN70O65GOK6UJbmfW5mDzz417ySM68iRnKYVlKxTimedR8m/jVqcEEPNsggzAQ3LXTzlgezctP22
XCDJu4amJJ6IjW0tkapOeLXDM+hR8NQp0PhPbYUcp7Q7flk0Gn+odlCgD9r78mKJK5n5BcJqDILo
81PH8JEbck5ZXhxXGJj15QifRC1N1GqSVl0R2Rtpi41HIB3191ifYGhDLTxrf6sj5mdMst4BsHjo
9Mdgb5AQfazDTsZp0IHJlPhLw1Zl/LN/mVQ8G+9c8fp3yHWZcjqEeiiv4qNRngJ7DBdqTrUhcAv2
u8zu9L6HFqvr7oqXA4nqKHxgqDsYMeChzWii7nGPVEObCdAkYJ1XnliQsj0OYIjn+0Hu0M052ROK
4wJHYZG7V3x/GLYpG0xc+5Qogi8GHA8dsPhx8ubN9XHXJ2Yq0QCrOi8eywr7ABea8txGI6dJT57n
JL08kp+Sx0KaB8O/VFGBzsN1CPzQiYkR9taEYj1igzZHqMoi/aA4dnu70c95y0OfBHctaitb5IqF
PQzddowW3Xto3oGy52Nj6AuxnvOTKFf53hdXXo5xlOnSLaUmbVv+wgq7UBT6NXJD96pLP5c1aDqz
Vbl3aCTA6eKrvaB/QY9TTQ5In5FpEOnTcai2AXpjfUem8Ac83cuXhFuivDwhKGiW3QbQDu2RMxQ7
AR5VQQFp7Xs+NFlXiGmJ91KHdjElSy+hyk7eNkmXipQ4s3n7A3Rkor2xPwxiBhXMdrPDT9QxOD/s
VbwzgRNoH152T/4bbmdfhZF/TEWMwxP9r3z5J4UWR1qP9fr4sLOUH9EMtNKrniE4HcsUH5uSpSC7
K+9DAZaB/M9fvAHQtvc2Tujr3yOGtdjppl0TW4MBFaj1d0y8tvw9qV2xbEGNyhSzl6I30pj0wEon
pFBmlYh7aIZkBGPTY5YdEt6m/s2RhsOFWLmOp9QjMWuaShr9wKU8mJpjg0F1+mCjZ4MQyqetpN9f
JzvlyhFvenYlJglmbcszB6oZmEr7/zGRVWj1Z8DvRx1LLpmfEg5NkJyPFDF3QR+KjJ5+REC5nIOP
0ttRNyE2Z/PwQTwDHi/NJuAwaDcMB3bOml2BzmLkg0TJhOevBuuVhTjX4iFyheDE9aDH2seoYzHw
+Xa7P1zkvp1p3uWkPBHSOgDfpQdnE21yPPWGpsOWAb9XbEkS3UPmXt44gR9V5yFXLfxczYC8Gfk9
5M0sD9iF/vwJoU2nH8mgrtEUOwUaMWeM8L2IwZl0wNkRfmTF4AcwxwWXn8Oyl7lF17IhkgaDUvNQ
KbyTlfx7PM+Ci8NqwdxPUGN+uEgH1IacqpwvbG/KGSySTlmPzJ2OnNW5YMlStEwhVt1XLYImqOhf
OjNeP5CTY01W4wJ8yeaCft6zXJyiqP/ok9Xxe/ka7O1ki2hCzp/js1AnAXw9FHF4DscbB2AgZPVs
chN8O36SdJghI27wBv18HWNMem758OAgOIkZD6P9wBr/NopInnyHneAPtH5BIlyDbFW2qN/dK2M5
G4pGRXaDhfI4CwL7DCc+BJJM4m/TKuLxfjWTiUsxpeMUyo4+qYbaD9HzEzW7jTLVFGUl6mhHgjPA
vLn3WzdA8/HiwYKy7fSmu8R69dsOcaP23soZ2+W1+ibQojMG/Kxno5zvhFfq2bx1Vt67rqdE/wUB
AV+f5YGyvqJdFF3xqs7eId6ijkzes6AG2ixYApN/wS+snEeSPOmr/wTlYxJQ04A/tt3xu7RxYrS0
M6n0QpZJ62DClW507jj9Nk4kePuohqBP1FxbF18H4okqOFESjR751WB1o7UsCZl3LSPEBw1q6EGn
9S+3IaGW5iA6mSzZAXoZK76EmC0ehEX9mYRGpfbtOyG38eA5L81p//SEXynLQqxx+m9jjg6bwfBF
bLtYXUXwLxoieXkdHD2cq8umND4Xv6M/Dr8+ccb6nl0cNeNVZje9Xhc/4lAyuHxOZ6PLWilr1x3N
tAtJKllu4w7KlzK1sYDcKk5w6jG/deG6ATa74umbUnZM7KY2Fscan04xioi0iOPoHfgi8/wsuwHA
JPVU5Mv7k0hZeIiKwcxGtu3Ex7brlKM6h83HE98v40H2C9Bb2YvR2JIfTWrHw7eRGkY1Mn1vFIhb
LAcMTEVIvM0YcVFHO+GO3cW/VMR6hu2nSAGqyS2P82747osM3vR/6cqM5gIT6h+0j4UvGqmGhvGI
FpmoSzgfa1/cORlm3jALLJdRENUHt3w0/xHbTsnfGrHwGk6Xk2zRcRqMutcOO7XdjcP+IYdovzvr
uDXnHoHSVkPfszIBm2SnyldtA7v0Co/yzAAIvKH+iOG7r2Ix/rUeM8E/cSXWiR4JYEv6S43kL00q
NV370uH2oCJOhJW8mVu98M1QWoHMDJPu3ZQyNhEICeb5IZFykpcj1Db5Yf+dUGUmq8msaAaVe1/q
Kmo99q6IDugpFALQfRi6X6TqlLKqSFNltIbz5I+tQ8AlErUwTSj76x6ZLOBydL3FPk9an3k8/QWE
CU5YtzfdP+Cxmt2E5q24xjzim/MXUAuTnBTuqBWMfAKSmXS6lXqfzafkXgO1eFxDDS/MqLaTIQ49
U9hXkob84mafLCD8zGfwyDFC26oJUW8xHmCeV5y4AzubVKkroC+LRZLKYkX0k/5gNamIfgSrZwUo
oWGize7ID96aW9StwohBJt2imyKy3TdQ5T93akBc0KxKdnD7iLqDolCtTxO2NspMA4Qa8Na+q1/W
o5qnAzbBlXSnScT9g7jgho0Nj/Noq+ojLAFJshi9P2jltJzSTvYHFFGn1nicjdnUY6FFsfDD88CO
UrIDRzMrjhc3CRDiFIw93icxSgAIrJUHSeewELeakeEybnVk5Njj37d4cNkkUwFKzYURVh/DCWa5
uiSrCIpANlL0pYJlSdLFmsuKR58+a20SKLQpzQRB6RXDlI6wyevF9JMWKZEXVW7Z7aBBleJmF4x2
6RkmGvDC1IUBgl8xOKV9K4wi5xDoPFU6O3kGLOmRLvwE/LXFD8o1fqdAzTwHQxIVyM0hvHQaBG2d
t8xQQWLtMo/L+SIOidWMjqNpjD5UIEvrw3sSj8OvnhmlUfjmfwFHWfuv/Xm+3CTxD1GMhi8jx4q1
PEkeK/PtHMEAKfolGE0cD8f4Jvq6sX59ClmFxBo4fc+3678MYmJIAg4ar+lxv5ANYi11VLI9NDOq
+25vsdZthBl+2BgCiWLfBVXDltbl1g9qyw7h2nEkYJy63DyAxK0wkiyf50PUjiDlX+16u86okW2F
2fb7LDmuVsYnoaUrtO00kt7SSlgW4xoqnt0wlkRr8UHn81PO9SYqIjkpGXggzERhnki6YUYNki5A
TunVwD5FTbumZ+u2Zj2Kob/HsI7Xdy/idHtrCDY1WuR8Ai6XvrVzW4xEzisWhVhuBr0kXgZi+dhn
OLm0yy4qNswK4wXpjng1lOF86YARzQKVIpYDRvGSNrZKWWC/HFeoqKJuNImUJjQstCfhuw9IINqg
yL/3c/P7CcWQAocoXruum5kLqa1gSQQYmf6jEzov82lmiSg2QiHaew/QdBZ06F8zVfbZkERPX/D2
wn/oxP5UkKM0t3X78CLK1UnJgiC30wtpnrwF/2G5EU85XrGHrDIMdedI9fdfkyYSpiizIxTnVyRK
rehNGv4EdieOA9rBIQSonWQ3lSrLxDj/euDR77zTEv/+GO+aovVZ1mljFbG4PRq+sr7cDW5/7mI+
dk77ep4DQh2F6Rd0JUfQoqy7Rank4I6LBubqkzkli/JJ9qQTnIqv53jNcoOxAIW3fAZnLIIqfqZt
3fhQH4blBAEOMRU2c6+ncNRtk5cSdm3+UTDexgLJ5dBWN8/BFmGv2kra75UYbs//OlEkLKVsVaSM
MuxI8i/1hCytVJ2/QBjRY1iP2P1q/45A8vxHDbttBuUoE/PVGvj3f6DxZOTJa/C7Z6MZYGnz/3FD
+0xrO5xgQVa0D2u/sTqFPndQ5iO4SOHifcOUgM2V9ZXtcuYstfYChguFV+0JHPCynTwixFaOhdf1
ohY0Vhjvb741Y5V2ghc3WNEhlhnsNFOjvw0PPk/v083kAFsz4MbqtT5mWUs8dRG0DwMt4l155vuu
x66SpOpFoiIkIijiTiTNYg7TSUyqXGfcXYZoqkZEl4Z9O6VxR1MAUYZrfp/kcmIfIBOUBkQ/tWBp
cj+a0rkvdXeo/uA/Vj7iUso6MYnfB3ADvN/ooC3iFheYBHhOk+NTvTsomqWi76SLKsBfiwYZtEt+
FHAGo8JHB4wsYYSYb+60lqi8HlYyjUndsCZuvsogM9AeXdHpAnq8ut7ldvwGm7xY5Ndhh+/LejAa
7AmAbLgGCbJRIRdEe7iGyU1zqUz5iOFP1vfu/M1UfY2BHngPNpzfkvITaSTKtQyDngz91WKIWfyM
uOaGGuccqsG4lxhChCOGJZ9yjG55ae0PVxHf5eySd+AVNIUqbZP3qA37weHEws5j2iuWrc62iMQm
mkd1IOBB3ZQqxp9202XaqmU2pO4/cDSRE2FO6T5bKiqfCBIqqFsKhNlSdSmQMjjEMSBQXOKrZfA9
4LCuAmmHk6hkibow5AxjIq4sTFhP+h4ZorATYzQaqxy0jYkvpfXR8DyNgBPI/LaIaXXRrhAmqlxv
uYSeeI8jREhDjMUNFOCM6xPoT5iZcgZU1bRnL2Nc1HKtStl6lO2KuZD9FoYxVlXr5OFkMW0XavsG
KXhRn0yWk61g85+j/syOSOI1eW7qExw5ZH5yFSHr7X99EOC4z5eavkaoVT5O8VgsUj3Gs5ecI167
4dl5p2tQGOo2Bfc5xxkM/CovCD+foOYAotz7IcqfNzHC9UbraMjEy5sx+ttGpc+eKwDHdYYb5HGJ
/f82hrB4DFjP9R7ilIfE3OO/3tzRIzf+eVzQlUFGkJQACZp8rnnlK9SnONTm3tKSY8/4qxHs8YWK
zfCyN9e7WwVtjzTqUBim4CnizW485BI5eB7nU5xF+vWIXub4PAq4xOZSAJITsyGCXwXqqbGW4/gS
v8vaL8WReeDK1sI5Zfs/cv3FPFfIC9dxLBMQlnylfmb77FYnrZScIU8ykJfRV5Dv1SzoPZFkMr7x
eqR1cOl6zw0PJZe7afWIinJei7qFOXSn2oAhI/U1XUx0QU0KG+8EUcRAivVuuvQ9v4gtulqtrLyr
wLWXi4JmFsA1yE+ksc+pw8+CgBWANSTri2bKtyX+hp0RRAap3+56cib5UgI0ybivLfK1f7+vEg+y
mGQ8GlNCfBKPbp0/TZWWG5K5RkXV7o6p6FiFNlD2TYojr8bU7SuGQfXGLYrMFwAdM+XHuWS+o58/
UIM1y+BN/0clKHcl1wtI7bI9vsSrynsDsaUYCSIOsnwVMPcGKAD21lzIF15+kKOcyATcsh6ZRkFx
Oe1YFzfjn5nLGEJ2vwY+bj8fBZYaXMeGvwE46gow5sVvOzDTPvkHdRNW1p0Q/4nVq44SiF20u3cA
0TnL+f6w9AXU1yatniEx7BUJ2x6KW3Jht/JPHmHnz5phtHo2h3oXpTWiN75woBIBEhH+/PhLnKmD
zoVSy5wkZgE8CthevnFu2wINJBujbO8YA+alYvVDd0Zi3qZGwlvDewj4YkahdRDDuW7BQHb6cW1P
4NE9pXuiKjBa6DXWWY4NfFLliXHDzdBfJlvejBehFGnSKFmAgeFQl7ji3+Mq1ot450wSPZJgwxG3
mmoPSiFLZQRnt1CwpnYh6kAe2U3sv4afnz/Bl9iiv8iCwu4o2bMTcocoI5Zss7f1ey1dhFy35ZH3
sVwRLj0I9JGeXJB686spA5klxsMfeKdxCDVHvQCbRN5NzRtJA5zvBBjwJWM8ryKTwKZ85Yr5N8Wx
OHuktiX5S/WKYKRSG38AqRmIaF0wmaj66lvcQ69cg+mh1thugg3XbDyLzvI600W96XXvS62SKc/t
uInCNt/7Zx6UIZfGve+XV5znc+Koejph8KIVTal4S+pAOj0Shv8jfHrHC2jx+LdMPM0BpipE4+KN
1WFySeQWeLGaqXxXqiH3zEbJTOweYRDK/dsFs4LkInNx2YKKB1yr8TD+AS15t28IMKtr0eDTTs4+
CqU2bFJZ8ADoM8ub+vNbzoB/vrXJLIumz3hFUrfPChxsyKYRbdFFpokYIEww+OGmuWBpu3p3Poy0
3fUTz6LutD9UigRsSYbjGXejAQovUDZK/buVfDiZCErddXducV5JDV5Zv2IVM7b67px0GVdkAThA
DmnsjqnVFgXEOoC0SlszgjslYZf/cklNsVv5LvLozxw6kFwwPLs1ZrGM+q+HgVxxZF/jD9CTA4u4
WB9o/BXExr1IcJS8u/EBho/Vu1DiOaelFqP7P0nqJofVOchlsLmrUvhfVdfvjoSxDg/jPtOgrBIr
nufksRuQU0uJApRXrVlNMpMOBLcZZMO0v6Gi5xdd2ER4OR1RxBRggXCU6FAgeBDmSaV9UsVuWkBU
ZC0ziB5VaXM9/ANeflvZ38ugHNSwuE/MRMeFoRZy1rFdnbQ+0YIK1992ZQU1c4TXhgxtj8UiakRa
0eilxFGe9M6AWE6gKkdRCEEmD+qEFzKeY9cRw6p2TC/XbnaTWYJDmk8oNZti5DRYXQQXEks801Wf
txVrBm2G8RZG+fu9bqqAJCuQ8RFCkRDTvYXYfct4qdgjLXstqU4PjLHo1WhVDGVFVXfacvWBnw6B
/aEz8xkcuGb1rThgrHgoXjCe7SgSEyenRHE4rvqRv8HVBJtJtBO3yTHcwsYDyIWFY4djtzaR1Y1G
NG68C0ZWYxkqwRl52/96BLR9Ni3egPioQ3Z/6Y+FD87vRvm8CwfkJI3M5jbMJ6VTlKqPutTcBNoC
qqTugQeYoNSrAZHSenWSgio1oXpO9hQep4Qk/ixHtvu+wnCGGqwD+wd51CZCrSxjlPkFjXuik87L
jTxwxRktvzK5XmCX12I7to32nHV4szEc9UADijGtCQFvc1hBVeODK8mEMmwn9GWTQkKIHpgBJhJl
qRlHoMKoUfKQlj0sApUkS5mlA7bLwEC5E0bcJxxyHCXrmCl6IIjhDbULRdHAs/eVBbNEqqXSInn4
ixKgGk8704VmBzzYe2ed81+ISvgLycYd5tfAgK9NTKZcGCFVr7xJF/SAxlR4b424QYDWPbQuL/Y/
jNzTfdeWoc2eUCDwGBi5iR6V54LYZNiI+whtxkgQRXqO+p5cfD0DfLC6466wRbpgyfy45kjquGqn
BaN7st/gheeKhke3h/qV+c5nPpTWMlc6Z9h5tTmbFhKgcJjnTy9usFASL1n5JJ5U92Y1vDO0jOFS
AUkhoPbC9/N3xk6B4mdZjLRmZQl/QsDSVsNHYOQ8q6cyKmAYOXM/tImbQx4WWZhHduW0lM3W/7E7
da3zCJVsvFegWIRbpH67sTrUm45mg15OG1xKLZTD6JdT/hohKpFcWd/gN7oDn0f3wngeUtJAOHCI
C9OnJKvEfdSAapE87ZBfmbuiVB/cc4qve2MkBpUBcTe524/cZFbcb1NL+GA4Q/JXQJg5J9gJmz+9
U3UYJpaxb6gzIm2t6sTMgWUVyBZvHCYfMIbG27es5QhVzptn9H96fhMiYgL8VLgFbKMafEx+cX13
3qLgV1Z9G6OALx3BcfsCSGoRRzcCU3bot76U/v8f48/wVVUk1dS9Z9CG0iCgaUsNwpdKkihdlj6Z
YgJ2VOw/RrB7tAYFR0PgP0nQQbnwXW38tltHMPHXEUJZQIrDzFYaDynqnxaPtqoXHKqtml74u4Fg
IFdM5u/ooDAsoZCVYFnLNOspxK/xKxTlxVfOYvlMP49hOSs40Kird5dtMzIJo7mGwLvWU29Zza4C
DYePzsquZ8cFkuYoczeBWy2o6RnPwMjgkE3f2hPhTG8jYNGoarwOwVgKcqzL+4lv3VAzGqT0Zn1v
py7xn74NwGI8IurVN9EcZQuiLU9mgS4emJmMPnIIMudyhDMXq3iuK2ZtwQyfELy2SHx5tNKl/3HY
n2KMjhzODTnvTCOulwUHjf0NlC53GpjSfKj2sCHlZTHMmqs7vDK0135DFaJlE1Dc7jHHBwqyBsZc
w/zOABZAA/cp58zX7JzbOa8H1d/zJEMHNyr9nOaSSWrh5eshC9MLmLc1LCdUw4+9j8rPkC2PiqBh
WpnKUv7OhjuvKC9Hg50/oMu4ZB6XHAxjf89h34vIpsE6uRkdx7HFgOOjWcLREpPZYZAJQonsgxVl
BjJr8SAZlrXxFxK9ixmZ9FD9SUhHXQ2TlH/k+grdhUjx2TKqNJnzIgSVcU4poEZa2FR8rZ7YfdRz
NWmWK4PNU990AsBNQOit+98Wagy9nAXyeTgThPKU+vLImr1ajdTJbYruL7yZQQJEmWDZDCvveiKY
CZh6Hlx/RIP9HIBY9/OyBkmpmwoyAx7v4Y6Rn06Dp4PgnFr64/54c8nQ+m7h8Gm1Ql9CvpaBynU5
6dCx3ZzAlZxtdW6+Ov5a7XCr0lzgbimj1aLgwMyppo9P2O0shzFUpw87n4kZDiDxmZBke9ZBPu0v
tWGVw3mnsHEb4Yw4rmlOBQM7s+c4u2sZEh+9gO68jwtgBt236zCLfZ4U5XjmKFZ9A+ehWYKh7ul1
IlNW/RIodB2Vzt8i3y1wH1RTsXjrlAVYP2mQdkyuKafVO5xzCf86MQnz0zyFZuFxu/0Oa0Kg3f+/
+0uMdA3wUyKtfnTPGcZHHKiz/5o7+JJFfLW1mjN+GHJmTI2VO2dIg9QNgnW0QquZ7bBgiFyTglJm
nBjtKC3y4stdgWdv9kcoFV8hj3vSevtyV77mH2iOSgW+EVjywz5waDqxA8aYv6It+unxAGZQxZv2
Zjq8Q6XwrA6CpSUl3tmvKPiTs7uXUbnht8yzwCe889xlPWXKoovFBE8tr7iAGo1Zo/O4RiA8OXHm
3GReQyXbbWuyAMsnH982TJZnK4/kO1+WosBFT/yA1V9S8ZB9vP8qvhmew3j9F2fOSWBNnV175Kd9
Dn8CQ7zbxnizBRQS5m0o/C9uIqrNxg6aig/cDvJe9xw4aDGOqLzJL6KyD4qYvDkl7kSwpYQHJILL
dnFdVCTsfgarpra4Ajtc9BwvAJjnLlCSHOBpB8GhTsTHsTIlSZ3CAWqjuS1b97Zpa4aLSVtAAWNU
0eV1OyuXS97vuZvvPxFRmDB7Xxnrwj0euAwjWAbSBJlsfI1v/w/CpScuDgYL5laxWTfHGu9do2Wl
127ub2ZJeZqVSQXkdUCUMuP5cxdGBh4JmJuLz6F1FE1kr5t2JA/dz4sIflCeR+uKGu6cEAupHzYp
cGEt40yQG+MlhpFoqGzHHcs84MrynYpkEgT3r55tyPH2ohDwRC/NEu0npsYBUZsQRStAr/PGSwIA
WzGMZrJGJ1YlyMib2FwCkrdc81IE2i1qefxeXY9Cz9Ajf/1jBPo6F43LCIx7q33FjWfcx/Q5+sJ4
NCtiOKPahtvE2K4cgoaPxyRsyypeSOYX4u3Rkj3aiTCiGEejiS0lhMnqLcVxBt/2K4HzJimfbsRW
6fTYLEgJHELoZYuvkl23wcwrwqJHtWtGmkWQN/J+Fqeg9OziyD14Kl/g3xNO6gIpjGMSnPCe5KNq
lAjOEyTsH+8OVpZNC+zBaWY+NmaKQWQYPJ4rZJXEQp3Leh8tjTZIYBv58a4iNNNCEEpuEA4S1LNc
kDTpWf3ve8tFnyLoGAsG0nvRYWuj/9wiObl+DhNvbPkd0u3/IvQHt0Bl6mQFAilcwBG636CYFjj3
2OKQeye8XqJZAqvWiyZ79ydz8dPvQksjDGBIqgVu3m2eCMS7QipCxweKvvi8wVCvU32Pkvg5V1Gh
fTED3SXkMiL8Qc3JABT27KlzLh1+ttNIjZJ/jzbKLVXnl6B3jFYbID/+ExnCnsUAT80RH0a92T70
tJmjIHvtHw/xFbAeWcUw7Cse+VQszkKy0ilfuNE2bB4PfmSTfN1nD9AGt+tsTu6A+bWDfuwJ1ICr
d8pR+2j/luaG6BBrePXueGDksFi2HC1n2sLo83fTZVyNjDWaeH917yL7niiKWAsXCpSW6k/Z/fgc
QQkgioysKjG5KBfcS75jJxPjLTNWT3oHYXsEAjFIZCpeuL9hA6MBsG2C4g85fL4fIYXr1pZL1XFJ
q6gw6DvQtFdJ8ZUdOfql6ciaMDVGNZlB7MzrlGZL7GyiVGdLjGuC9w4k4ssVFvZaL0qOVAYs8v2J
y7S/E5h2XTCljHmHkMhWpCWwU0biA8BR3/eLR/XThcOO/LVwbfo+g0H1G3gDmPvMjj3eWeV8iZcA
9NVbfVLY5knFw3zUY1jS7h8snJFnlyta8uDSZv02iv92fexbBEdIOrmaQg7ntla7QYm79hNVqXkT
3SPCXg5DT8e/6ojUvfpFZ85bjz0T5dzteNSnIVkQp0IJZzcuYEyO81QV8ozCnLBWHxIw/0yusoML
yj4I8ecvb0h2abXYvCQM9cfSyMKfB4GYbo9ypLlxxDhyUufHw8Pd8J9WZY6S8g7k6TERI8f3bh1k
Sn3lJyiWHCImEcyQ1j+qbMKgJOWbUxc/SRgu5UWrucAcNMfMtJ4fArF9SyoYC5kFv7D+xg7yvbK5
4ASNoPh0YiFlzdQF+Y81x2+N8Kl9aS8N3C+3K1c1UFjZzyQvBbODCeSOtg98/w7G3nn9yF5es2av
FEEKmxYQf2mv4PZmvVMM7U80WxkUzA/WiELpdEtONFKCf3AIuSO77eZn9c4fR/agUAlxSpiTrcOS
Ims00gjRGaCJ7Q0vfJeu4n4VBsBF47jksdM5+XFmmfJ8G5fK2DcVN9J99oiOBiSn41SDjmAGW9fQ
4DdGAOCYc1/eiGqVIsNdokh8AjFHs9Ju2HYS7omf7fo99RUN4qpBj+Fp6c/z0ZaNwJG1QbJyF1Ic
y9bmKDLTDEJXlgEu24M0N9b871uMTNUaOTewglQ8m1rcBmXbQY9TaTGfpxYYKK0XhgXbanwGEfQb
OfJXbH/TCbWEz1zI0xYvQBn3OYrJbZeM5UNLA1fISwtSSNwrVo6UAUDXMTFYdU+2xI0Po+qhaiZ4
kIhhdZdFWxBd8P/pGeqwazulDrwE0WtC6T359706lq6570DBgU24HGDWO+wmpOcybmm3+2whHZo3
KawEpFaHiwEm+YFJyb7smBjBTwlhfx6glyc4LJAHoTxGJ7hJe8YeV3Bh5pmo3M2iqrosf/pyb6jq
HHB+uLW6HaTxaAAhmBefciZqXgHFO0p4Qe8mg1xzHkJU4ql3/tvHJieiKHd/VTobSrB2TGWpy8Xa
ql3G/T/4+/dRrtDugHJ15gmuJW4CYvZTR41SQKLXtKf0K23/pewAJRfZkFm3c6+SCmmidQaxOhOS
ascDllFMXSqsu2mmQRa27ymOnp3Uh643RmZboVW3B/FtVwONPw2jTOQRznfsnJ8wPiZRNt6Vfsrv
4dKCE5wT2ejwQNC2kFl4EDfQ1ZVa4xZ+H1nlmwyU0ngtTMwJoYPTSSAoYsxsunYxZ1yzdpTyGLen
4LrbMndFWYQFHpoGCWc/pvMhwdFeyHT+c0SoWUjLXfrF/f1WDzhCGJc6SvFIdHgSw+bQXkBfJpdI
c2auirLVEZp6ljCVAa7cBDVRImkKtpENxVLg+3EnKc+CZElsNChi4pDkH294dMu4/PCYNQHs/ERA
roIs6i1Y3l+r60zAEqBl5lr6UtX/2GpDvjTUFaIHfD6keJF4fhXZfvKKZuH97hdDPxO3ZRxmnQkK
cs4I4ydj3OiMgxPI5fS+xyUkV7rDe2n2ai6o++lSumwQJFJ6UsRoz7s+KsiwwkfPVLoOAhS9ap3T
bdFbfc+KW06krzjzkmYq11xdOFHNmrqwNnOkS2VRPrpr9BNRMSc99ZRWNjzVy+GZb11OLZICPx/a
pw6U/zzjMbVKlWoGT0qRfA6uzLk0zHaXOtDJ3tBVLcnGiLdMiOxu7uxbuquVMcEzxSPhmXGu8AWZ
sK1NG0w/gaTBkqPYxYeUL5/Zi/Z4cM+4h6eQQqBWww4DqDZE/UVY1Byd4CJ4JiiYHI/AinGv4VuA
EGReljVsZXcZqD32h7nujAUX9OfVakKxfEWs1c9BT08jF7TXcCml3YIfnavvSWpTnU+ITc4gxhhH
JUwNDJVR0QP7rbqmLagf4ILkt9O8os0R5JOmLiVGshbsCg4FvhhFHj5goY5HLcFjXeKv0HOjxj3F
FEtcMxHL+BrNlcdZ6AmOFw7uHzDaNdH0PTTfu5ST6Vk9DoGRtCPDfl3LGpT3UZ1BRDuPtWYhvkgh
9MESYQ4xcGJpogd5CSY80rJnfTBUoZKT4Mg9TnOttvAkExY/mzApVNa18tNrpCpqMyv7+Rs3d08s
NjUtvxAKw3DFNl9dYJb2WXBfd0lTJPczuRBGDmbF1ZdSghgd/miKsxaQETwDsaGxCXuX+B6RWP9x
VJN1k+Hh/6LNeKuabYZDgrKxICj4EpZUPKOx8WWooC7HI9bbAL+tjYMoQ8uUFqig+HTC09Z0ikA6
udLNtaEgGszUZfRlQvP0bfF3CXgovS0oJU1mXMuIN70RXPL6h0rOUpJ8jcfECEOgdbOVgBFNDrzl
2QSiXehtTQJ4VywehJYSXIZgcJhddxtPikDjSJ129PU4xWuG5zij59De1yOJhWwr8lGCmGmMKrKV
vYrFnpKIyKCq653Em/eIclG4Ipc8VQC7V1BuHWq76+1DwJQU96l84dmbkcv49Mh7CojjzP+w/HfH
UF28rMFDCPWSdpmRX+jINTCJPp8HOu06/XUXjotEOi+kq8z/Zr0hbeUkhfcDzJRZzz913qBpxSOK
FWo08L7X9bGQo1JqbF848qUOfHypY0Q98Aa9aeV2lRLuTKRYvZJ5a9w4TJtlYqG1dCcfQD3/iFhP
LhpZLICprK56HvpUdfcNcoVu7pThfs9b8z5xwI7v276ivEz6N9Y7Uh+v40lfXXiDFy9m1X12n+GW
/k3IrPrp7FSZ1JCarEwg+2UDzB0fUt9BoZGVTwSAKs1bC6aG4/bS2hw3fEmBMDtcjqoHU/Tp1887
inn/3qoHVQLgUdkxxy+fyAwJshRUpnV/N3KhTmsgdlglS+nSD2XH72IlwERKk4rXvJpz/QDxW25b
YUgv85jrHOIPaqZhtiqivmaEQi0SH77T42BEmgfKSITKy7fK1noWtoAfDgVVVXRfUt8NreDEG61T
uinlqwzxCAeZSL1D0poXkAPoSWFhwBzJjYGpcRcUjJbCZe5Jvpu/iyCXXLlvrGzfeN2Wc3MCiZ9w
sp4lYoeGSnQ8Oa4RTrcq7CZfcPeun7y1wACdfA7mFOSBNyBYXXh58DdhA4IuR5T6R+fHnWRG0Ynl
RVNzE+XYwRldqPcfMHgUIobKkq5dMTqxAAA2BN9Z7arjwzRi2dkxNc3yMnoyO/ybKmgmpQJOO2Ui
PILeWbiuzGf6Kqq/NxmrVLapF/hCWv4Gy2rROV5ZVFN/PmGyQslBzJwxPDIG+z1SCYQ4hVD+Qs4d
SOJ4HXtUOrK99ff2t7zofi1xmLRj5Rph+wtm9BM669Btlvqwxvici0RQDufCq6IVRw+gBnO+wugF
xSy9fX5tSXArugAGTNU/XoTO1/244IdsT17d9y7TJeQdjumc+DIGhcV6mK/ZP+LwhZ7saAUMH15t
K1Q77a2TEQHNkmWWZezzG3Ew5bRp6OF1scmdYY72Q/GpoLvc9S4P3QlZEqC4m0B204BDU0+za0hx
gNyerVX+BPWW3x8YvEDfupnrflWJYkE4ziXeABRgnagUKAakMVCfimH1f6x+49WO7PwsYLxylXNR
zdIQq/MBxIpeRO5rtXNSL9VL0uIm07Ougveact/iLvOSlFa3ilZMfUkCUwawEnOKu6oPbkmMz1KG
TufSRDp8Hf3YoMGE6tZn3HcBvIrZVWmdyDpe7IIi4VEQgbBTHVvMORSU00fFcRS3hAA8Gfp6yQ9Z
jF0WwisJcP2pV2gNQ5ovjN4e7RncQHvVCck/zo8/B7y16JtCXfpHOylB5b19d0ZScvS8gwYbN/jU
5LtvIArwisAOo6dJhEzeASH2QuGbJrHf47924LCOUv5/u82/XkVUR2sRRfgY711NSnea77/i0nPv
t4t4FYTsh56Uniesw+Gg1lB8W/P/XZJcnwBfgPp7W6GcJF5syjA0azW2dFaF/9Os8tIJPaYcC9u1
JK016jxOlmQV1QeTvY33KOkq3Rwd1KA27wdev2cabRINtrVPO05XquMUAD5WXF0UWU0WBAho7w46
fNglYqQ51bnshaZKqAhBAQ7ozKBQbKm8P8p5W36wJ2K1T+2K5j6BF+R5bphe3gsCsxQZJRoMrLz/
Hoz5bmPC0/ZmkWdKn/58DjSy8yT2IvNap37g5a6MQ6SKd+66Ua4tfloNRjtjhj7/9HSOn6A1E+bK
I8/wSA/1bbiu0lWIisNl1WDYPMCvvIgvaWgFU9fpFfV+xTTYaxWxn2F8JyK9HAX1oMPCrc6PwEGg
Pjb6roFFkA5kLlATG6mOZ5TO3Tpsm9ByBOEocZ/j5cX/imYLWqtoaJknPmEHQtSi0pVd68dPfWqw
Lz5aOdCS/9n1kTuutEWc4QeeDDeZ3/GsmRzJHvO/Xf/uuFGIuEKKNhb6J0x4zQuHZCyDYF2a0F2m
WM3qwHLXzqkHlw4JSPG8HrFPm1ZDIvgszqI9PqAmpKusrk36QyZoZpN6XnW2YzrYJ2GD0VW2kOu+
zmnYCjfIFEBvDyov4jNsezNRfPujc6Hargg4wjTe42mwnvJsmDw6xjRSp5ZEXu/tuIjUslT4NiGF
lU8jqfns7vrWpgX4ckInhUj0T8iXvjYJ5ECgsWhSPAnPOwWM1YBicvwH1m9MrUpMG2R/VXC66/od
+fEVYXf193DXYbG3pADfnDVe8vGM3Sou9RJDHahC4t2CVf0EbKUTWarpVybjQ03JNv+ushtQ0H3/
L2uXYZrZMFJBw929JcNuonr2xU+o1+b/sA7QuKE/A5ulEaF14HSjz6NzQfDPauhybtJ9PSFZBwNK
k3l1oYXnpVb+s11ReHfl5PRy8/cBh0lPKIHbos0+yzL7uI66kdlsOPzg2AlGjBdqEkBz59qoXdAS
1jU9CYdzRSjvP4i3usajhNjgtlpoI7JU6vMWFbYnjifaejLhEW9KFP/yIEJSh//CWiutuEsmVAY2
snz54hPYiK+Tb3r/29ufXd3AitcJvy6aKjLcJMaB6omibqeLtrPPTTuE+oJIJ4EnOopKchtB76pY
S1NugzjZTdY1FHujMcwTUW+iH9f7RJcMRi86QKtioLJ9EfhdLhG3tVrEcqIuXhUJe4g15vWQpzE2
nPwGko7Vj1P856CvfS5zSl82VhkYNCZr5FH+P4prKWYIrfp8w76/cZuMwGfwuRvv+znM/R36Ho+n
h/4qFCI=
`protect end_protected
