`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FRAqbf+bBhoBolBVK6TrIwKUW78DsSsfBWjtXj1JPdvxkcM3LCcmPeezeH6aX5QtTzsUbG9bCs2I
lmUaopyRUw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MjXI3IjLE4KlwEz8vfshwXOe4b2NF51CKCFgNzY0hEwUT7k7DO+nrfwJFiIXVpgPdo/Oawnfdi/8
0CG93IispXEdzpZOCtRdNhlCpt4R6N2539jOse5/hR6nmxoyFos9nUGrv/lZvOieg2BFwFg62UJT
Hpbop6veymLH+ejHANE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i+vKqME6Bey4dIN6F5CPdQbqLcImkxQ95oyV5SxgLiyrnuE6AM60BKb6Y5qYdO4RDTWcko9bRNXA
yV9VCH9S5+iM9msyn+1tw3pwZLbWr/o8ilXRd/oZ76piXgyqn185SDG2PQ8UhjnECD7wufs+5yIV
gRJEAcXzrOxrokorXYfhpdhxfI1EziqtCl0NNw51It/YfWFWZH6l52OBjEU8g0sRpo6cdPSp0+r5
xmAJIBpa72sCE2UMsJMv2iE6fJJsGQN2kmKvq1+uhlBWcdm4hsPngsh3zg2A0eQL+xOweGrB0ov6
27mLaJUPAsZIutYmL3jxfE1caX6xWuTnPKbXvw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
N5EqB/pvpmFhp+8QAg6OdM9dZgbPT4JrzkHAeYIIOtzb9dh79xG5L9w908aLPGhdHK9mThnBalFw
mD1k9BKFOKAITZx5qU6oaUiIkp/shLqWJQvACL3o0lmplIp7rHzdz0idCrxUls2rXL9MlfcUNisQ
3XptfiVaEzgAO2qiE25LbzNYI05ys1dpNsJPeoCBdgo8/D3Ma68ajgOuulyoos9jYtdBYB2d4k2Y
cKRer6zZR4PSiU+s9VIiKNQ/QP5B1QrbdJN99lWuBSsl68NMPXkm8xGLL1DLbtqOUOTRgGZqOIsB
jqIsB6GOPb8dIqIYzOxNZCrucrJnVF1b91GDKg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t8nCUnMrKJ3EJgrCp6NRtzVYvbxHoD6HUbZONVvgxyICGzjN10XQ+3rP09LrJ2pBJA//1iV8sADj
NaGf1saw47eh2JTlfEh1laaEvxg8bDNsrp+YdUgHpoH64pVaAzYzLNcpfPgt0EMCaOFivCTxc/YC
ggtRPQOHh1mswdwrtQQ35AgNVwlBFLnlRqRPyjFGYrdNJi0AEt4hbbWl0PYTEiKugnaZGhiMXWcV
Pcvupg12mIVv0MDZSoltbeatNgH3D6uaWYFDVq+baMnbPLW/6yXoInDtyYsSuE+bZ2oVW3yrv/tZ
DGAPNzQwOWR2uXcQ11DSDJbuIf2NPscYQZdwnw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D6r4Z3T7oUmp9p00yfD5JmIkR65ntr/QzQd/90PcfPyw1EJx2355cx36goDZE5UcMBzH8zXE1G7V
WnWgFT/rrLyFfGQMRun39Cr0o0pnRQ2Hp2iP5z08FyrZGyus/dREHDrILjAhPt93glTutktc8Wrm
QSUyRcwb/l9ndDuIaVQ=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cvz5zjvCBO1FAwnhtcCOzmVGagQGz9MZ1UpzGL8icgDrfTtF2kbD9XarAy21MMSGoFzM3rmbemy0
8kkyfqM6m6xriamxYCee9J/5m3MPK93kZ4JB4U2D7pRzyQNZKhoxjP6phtL60r0rpjGlMV7LPqGS
SBin9W7VChH0itaVRnaHiK3SlwnurVuEY/DzBo2jT8L/oqnsOD8kUTBvoc8+nA4iKuLW/R7Kn0Rz
/UZPCv48/fSv8RTZM+LS2jPkCSDokLQO5ugyvU/nYH7+RhPpYBAE5+wsjC8eqZIV8EawcQRFATdX
VKdFEAWt2dGQFUdnamBkV7SKfgO1Z2kQouVQNg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 565792)
`protect data_block
foAKgekoOEJ4soQ6VoTglWwIosMpkVsvulvMziirZkEPVYjYJ6NtiA9LStBf1uVfNZTcZRaStGNf
1PoLih6jEM/0mK0mIXhJ6kJYLMZBbx/YqmQtJYsV3jakUsvm1E8F+LJXlRH4EPO4/dl4C7nxIXPD
pVqHxSK0zXmu1qOvuhSBt3WY8UTQ8CcXrhRmvS2E9I0Kh7JF9NXQxUcyg+xRgGF/Mn6JSEoVFIve
GupZjkTDwi7YsWSxfBLmqz35oCk+bTWQWTsDMWqxOvEIYKmDq8qB8AE3EXMH6Wd4r23E4HQXct98
U8ya1jwuQHGTswXegaVmmzQvGVc2+4WU5QJk8HeCyvY/pmnrgwrmoEFEG5K/2/9kBjnyjbuIW24V
goP4C1MtOxFwejAl3aKkzDiyUZnwX0fgbGYM56L+P7F6q4AHMksm141E+tiVp9IVRLxFmO6Ilc5+
rM6fVqmvVJLqlxdKUUyosQn9V/BeIysdK0OEq3R4azb44hemM8Tx4DCzMRqz3pOEWdgO1BPE2uaz
5Ti0q8KnKiTAUcAf0l3zsnnGO8SdF6bYcirkTHJghHKUglj9sXgtADUpKxfKxeg5m/Gypx+QTFHh
SvTVlFhE05DRrsVYWr+3CtzEfI4NCjy8ANey7orRckGrFsUqNtHlhtRguwJYs6nkby65cN47uWl9
E1y+VsKE+7lZICOIEMGdwVMpHMCQ+FaNZblWOGTvLk98ZEwTw5D8FVIsTxJF0sePudCjAetMQbyL
PLBSJ/5NH6vvA1JGvm+f15TucE+pXozTEbiIFipcVttTX4x4/bbmbPqdqWn991ySyxcHsr8AhfZl
ZQqGoFfcHmKwlHG2eeXsndt7qEO0yk2UXLvGV2wS3OQreE8mYZEpor542EulQ2f0m95ch8MX/Wto
SadP5VEK7y9MH+yRHAO89jJ4SePmYm8d5tPnJidOVcenxOF2ivAK9gbiNs3ECMU/MjwB0jASxLui
/mJuqTIhO0ULtazKaAYK4wLBdsZDTD5826RhEkzuRdNEkCA8qiRxGYY+0CNz8MO5EG/EVf/vfAZU
QGa4O/+z/DdzPOKbxrvMFV8yXVc41oL3hWFLZo4aL+MLzlhpPts+EmJt+xZZD+gvARXhuRRk8U3T
/MiKBEEGr2fQMx0iIWwwgisLGa8UkAF4d21fdXviDz6IlIaenPVP/os2Ip6gNCqSQ+gUmUfvNTiC
uB6ah0QQfMWJnh8N8UsInYuatiBGXZdLiNkZIMuY2mx3lZ/zlQCOT/ClnPFXvNLtRXO8ljnCQJxD
79Kgmtc/49+zqejOKDT2CARi6eVeeAIBFZT33svMNy9d7QrOkHFTM3tJgtdAI88XezVlHYP+kaLy
hM18qez2KkmO92Yre56EtI4yseNpzuvLxwKnrI/4e9lpVQflnamxl4hDO319Abyji56/XaHV6p5u
1IlY+3wMnOUthTReboDJkAajiM15HBUDatMImApNq9++DO3wDY0v9AuxAzxF8YTOHil/c85U2uc8
Y39XBrXGmV1pc69WXZekRJ9P52CEtkMqKIby8YvVvkXGkWcMnybkGIKvgXCDkiBd0qOMUKI5jvVy
qVXnht7tpIBNlM64syfo8qydy3xHtl0sUHpxzpG393A0q7UgWTDs83lns6v4jnUjT2BLWP8TBps6
x4JWYqDUnSwLl0jt0ovgraox8vsoI5ePZlSsSNwtM1eAgpXnVI9kXK9l69QKjtTTL8kZbiSZpgZV
MMKjvvOxv9tZutzEE0fyEofc03X2MmQU1tzlnMBcKcd5pWcpsXaEhFoq+IdSqPCCptgJGxrSCa9x
hOkL9Y4IfoRa8gTK+TDmRNx942VdTszQqAafiOkPsctFfVd1MBgXJVNskyKAjc+9HZqDkcTjjetV
GPxsdJdu8TN19Y3/Rl/c4GBIW4dmp/fs07ErZ+v80FA5zAUpndAf5zR0bHW+QgA8gzzWrhMhfvH1
2kTjhUC0ceTHwTCqdAowK2cRJ9t3dW6R6g7V+37m8FV/LBuQA1Vl3CF+LiQgI3gC5ZQ1ko5Zj3mS
pTjzBUbumQ2gIkEAW9QzBZcl0/oqN0qd3b8VGRmTQHhTPAqmRj694j/8LQFvwhbUebqIgNLPEzZI
08sRUob558il/jF+yrJPRKECU018v/O8EDbPo5dCjr2FrtdPSczH/mK93QbT8Oz8Y4D+BAiNN3k0
IUYi1uKlACWQUNRJqh1Y7aZkZZ3qQx4NXIE7gHju9fFplcl7S9IPcR1gMxZAvEFh/sHwsGrN4rjW
TkuTcCaEyka5IBOlznLANZIwLxwqwgTJ7L91wkPDteZTvy1rpascXlOILRdX8Ee/1dINF4hAV17p
IIVtzIBLb5IT96ktG+xVTF7JGNEC8JWuPfCsq13G0p+3NjlPwRj88lxhw4od0OODHSL4sc80JTU2
A5TGiZu3UC/8P6hG2K1emEhRWAczpABez+kLhrPZdrbz5On5ULCUin+fNjtj+R6c4QkQ7WsoJ7/g
y7moEny5cYlpfjvFF9yWFBMAIQ991eC+PQRfa3eGuAj7o4l2dVYsY81dmjTzMVH3JD/65bw5vkgX
uAR9DFj5DvtPNRTGrqg1uUwVt+ryG97wI+gxzr0Ccicqz9z/q50aYxbnsRlt1kJcvJ25xGFRIymQ
YVWfpUHhQrPwaG5u4CkhLYRDLLE0Gf/RmiImSpvACYL39SH1gVDtxXIxvQws3UNQlji4BDhU9jiH
brBrjK54l6UvkSlFjGj0cHwZbuiWXaVvXQNAXMOk7U6mw7Wvny/ysK/NzpVQzDWGxbwUtU2bq8Hz
loLvsy1j4gSBhuEgORvlDo0NAPwJZh7XNazxKNTCQo6NwOfPjqcHa5O1v0DcbnF2qQkXrT2W0Tss
TgVuJlDWhqAkZfdeaGTJRMTR4R2/0tBpuIn9TJ4HtRSxds7hsjFqR3oA3IUAB/Zjhaz4co/VKzJN
be/9iVN3c2wqPEQzcv2z6s0hPDaLw8x/xv2D9a95qWMtUUXBXZ89FEZtD4L+SzQxWvX4ehfzgR0d
qhH1AS3LTQ3a/Hqo1NgVPPxpkdEX/JGyCwcafmVSwtaLAyIvpJnD8U1OnKJw5+nt/zXTaueesNsy
PehGJ1/geYIXlONp4LR4gxySBql1cBiKIbc+jXXB03LpJDIi719yE1eH6Py/GlDKZS3ypCK8w1c+
h1qK8/7YbofEFyScSCi4XtxFEqp2iCq5kgEKYJyl60QzPXCB1bnGQvKpq2Nxu61tk6n7W4nDDoCO
sg1hLcsB7G4aSP3nyHddd2NqSrPdUIrB0FwouhZKl/DQ2Y43dy7sDZHYlH78zcfgftJqwas6Vm1/
0CkgionzNzuHH/vf7fP1u8ADr7SXPsMvVmLbIp8U4OT+sEUifUlKERXHBQizWHIaR/vbBB8eA5Sl
Z+Neg/rN5SmMl4LmtJIVQmvl4O6QENuxOiXoli+xm0xXGkVWIyrpzZlin0oQcwuAIrC6uq17s+vh
QJ/yl20hJPnOXnoO9JPXhnY1Jke7H/XFDSfdPpBb0VfH1z49xqlTOT9kJp+Yi5td2D3OH5EQ7ua0
Qq0jffvIUedmDKqvaqtM72hJlFnhHAJxQuMjGY8LB4uI6QKqaHq85XRRN7vD/tjY3ivS345hkJRB
l6XXaLhbNOiiFWa2e91Xi2AnLjKQEVi0++nNnB7a4obGQxgLKrtG1s+DppNz6WHqIX6HanlPz4wf
IvQBo+Z/O8ppbybKdFCvivy2jc8BBQaKjLsn+oQiFdVfhTOQZksTnVT/l/RLhMTS382z0xoTJHoy
+vzCYrQrD3+LREvVlxwkUlNNK9/xoroDikK5Va33j6/at5UOnq3tsM4lUCx+NfPJ8op8xlm4uBRG
bdrU9EcI7StIojh1vCZpNTZytAeI0DdvRYq7v8AAudKKeD79la1L4hpOnLm9EqI5IE5jDwYOGPPh
tS1rmfAOe7NV0eMTeLlKHj+9Whudpqmo/Z3lywaGjm62G1t2ROdmPapg/y3XRG7fNaSrKsr69iUt
MuxwipkR3/7AfvEUif+pIGyhs8AJbJVVgO+jzyZxHSaF2u+SZZUwG/SAE+GDZkbBNHkKWBc6iLCp
KGpFQ+Fb1hylH9lfdp32Z0vUcwwdkiGZzJ6BEJqXMxpRfSK5CzB/L59+jUknlRcw13Ra8dPyG9Po
GPuxLIeT5Oex6qcAZIJ7Rb2GrDHBAxYjpNawRLyjddnAGyAvC++fDn6u0qwMKbX7J8dP6s4H3CnE
7Da275lC8q18R83OCm5uJTAJEkJv8AZG5zfH3VfC+HixF/zWOqJr25//U+EakMAAxBftQ/hjup50
oIPgbtoB/iplxB8xgrwqYiOpPxVIVtWYbYtjU8NtRxJd1oXJEY0NNyVVqcPjtGotSAYnttJgSNnP
Ox/M1fbgY2Q4GoIKNDjL4iiH30a++ql/V6lCc1BL2N+aTsy0lPS7ugE8RboJ9Hax25whnwr29eMz
Ha7VhI0DNkMlaMe3WaozI4vW5FS3T50iY8JW0g9H5DWl0jc1qcB1r14kZY1FO1MW8TVSocCN4ln4
MUdl0uNxb2FJ6dc3p1Xv+VCxlXaOsLoxsb0Jos4qyLJydS4A5z48H6aq170fixs0rXGXhxNzztnp
aL84xu36gMxZytVMuwgOT146vqFzAJehX+3zPNjZeXHWLA4iMhE/7ks1meNRo+M03vTTLV/g4NMD
cOOl+a3NsNAXAz8Ji8fq1NieQt7PkgT/RMsnckyT2HcdwnjLztZLYb9GVr/VN43kYt4WCAbqf9B0
V7BHZJjji9Nnm9R0f022DC2ctRuSpA5OcY7N+x4Ob+83mrixYvVHyDSOExKTc6KZT9/rB7QmCa9H
rHCc1L6eiLWutk2OzDsp/SuzLsI4QwFr1IO/2jwbNDu1qnrudSUcR+C4+Pl1yBFBmycajKOAkHK1
4cvvbGuZY5JhItjztXDCezHpq0kGtUrpZKvPUmJMynZ913dAdQxjfmdIQWrVkSEWsDbhKeaVDR6E
Iohq+CGaTZU4VDvL6gtm/1S2dg6dvmWlYAuH802n6BE+0nrfqCVRFX/6lmCzcXJZwqBSlAyYwDw9
r0XY4zNYSmnI23KhtT9AgJybsceSvyl1Jc+gABkJv8gTEAnV3xNNoUxSNF78RunSYtNzSF7GbEN0
rQhfvntKkYf8D2YHH/PWvOhaQ/bbU/IhbcO1iK45spsjT1W//AgDeoL8FRzEW7oUat5k/Dm5WtUY
nsMy/OdWVwqKjSBjMGg9yE4neqcZkCB+olI8MJgza6z1lFOXU71Qiv4HDm3aWQEciIhKiw3fMzLH
DjHqSmzLE3/QpjstU1IbkW8BqD9TdzSk7a8KSjoCwkdd13IlEWzy4bLEwINMg6WCfQCvyg8qyQJa
zFrQWzD+Xbl/WWHnwVU4p4lzvp6J4TBGOAsHh0ybW/mOz291GdNu74uMSgNFRJsvtvolGQ7oduMh
ChPLQqz5SOYMjbP36Oc9Wahw/eQJe2gBX9FB3CNFVqUuASQICYCntiAcMCznfgm3ErPYiQBGEw+a
j4q/m6H1VhveNGmj6QKem0uGgwoxKHGwcxWFgjySvLKyEON3hirvyZnXU4msMXvgL6+4IdNh+jhB
rNICc3soZ69Jmg6WlEOIXFGiba0GfrtlwByQGsTzAV/Sodv9LPtYoMwgcxDrV+IiT4BbcecegTcE
3+4CJWJTJDmLvd3ITHD0+dNNSrO/NEcgl1Bz6KkbJ9Dgyt7tiwBMQLECM7gvOqr3WjakrYBEyuKI
PDxz0eueFcovVMFetua3DNK4dnHok5IxWNlwnppTxq8floxuqr+LAMKj146lrXkz4ZeM1S9LO+34
/LE/Jg0waKlhwJ3QEBmCgsnxuLNIGqvPfuVxIrXIA27TgxBlGA3IEGft8COdzitHsVmWYbNk7ReF
kcZMdWQ918Xjqu47KEaepeqm76rJ+xi0c+OCWOlhCecUhb/AKvoNryDgnyVEdCnX7Z8at/CLagea
nYB/gU17hmMhdR2biVftiSSaZlAUbENh2SvFxoztcjYAMeTSJJ1quLtJnYLFxDD9oh5WAtHDSc3w
2SkoJFoiTQguyZF9imAd0cw/PNfGRlfEMGjQpzOxR9U1E+bGCPEXnra8Xj1zA5Sh3JpToFXwzwut
Nkna/W8VNmB4+FCgLekMuFhd1joNwJIuwKIF51FgZpe+Ha5NVe2yfdofkMfnnhWLoDZwdR4La+Fl
Vv37Sa3AUrsVqI+bMytBoYjYu9Um04Vss77/ua1gRnG8EJLeMXCOBpHR876FXiyiXC/JgAE02uGJ
nQ6rwCTiM8pPd2y257t9ZEvEPjsbcHot/zL8i94I+JxVz6MbERqujyCaiMcEjMXJyy4JO2NRwanu
Kj3JfoU5O+Za7O1+BrLtRg1ffBA25n2dEsarkEob0Ml9qJXtrJA0l6I5uynLBAO0ojerhWwoZg/H
vcJuBxFrbe3bkOIrhlygj3nNFb3/5ua+RwCHxkCLXoTG/IajhKBytrRskzD8s8dWlPPn6pQuieeD
gYTKyXDJ3s7d2KT1QkwCNpIVxUp5t1++o+sY+qDxLMZz3KytIvdRGXUqabjeTdDNxgldjeXukDeg
c/L2YIXEdIzPS52dpw/rJCLo9R0T0fLkZxma1Mnadj8C6sK3w235nYQMATpMB6fGXAKZcyY6uJCa
aJ4O5n8qG3GR63soQYW+fb4Hlo83EM29KuzEZsCtq7NAxdZTrglXS6UBW8LcgceGYbBPSnBulbv+
DQMmXorZKKcD3pWWJR9RsOF7Gc+OR8AmGkQgUmsCa5V3nU2OCZlNgxl8x8C+7/fSoU1RpbpXCeAe
nXkYKeX+SJq00m75XbP9T/cyQDtiEL8Fe/E6gjxQ4tYdWXHV2ylI7kMOISjd02KMJVWDxBz/10r4
FGLgiM07p85bWIfqCUo+Rqkb/VG/sYdgCpw9uVouV5ueAXNEcmXGdYbSrYWEb4mtdiR6zNhsbf0P
SZ1Rnj2KSH//OHJ2q25ompwAdEIi2wE7puqkl5mUmm23Npx4RrSQ4V91s8vrX45qh2BJI51yEeD3
hVatbrXdv8T09+maGN27OYE1NU4mZn1PSXH1NjV4JoOqO/nIQfa3lwu8lCjmwId9M9tkoG1aBx55
dYe6KuPIsVu4NsYNQ5I4sPns7PjwF5yfwv/X8dX+6s5gt/8rKwy3pl4rZduMMH4n7/e4+ojg6Fik
Fjo6vALJkmOTMcYwYeA5/MkyUKaP69ZIQpNDXPwyK51Pa8E+brX2b2YtGtFhIklSSVs0VHF8pc7D
VZD+qD0jZ8UsmpGGabJ/uvds1zN+yrvebs8sXaVDwy405pcKkoOKFr8V2SrN5QUmnDwOmBgXEMXe
6wqp7CTLxuPU0Vf5BHokCzb18f6Fd1kpVufzzFyciwDca1WIjmEBlbHKQRMSniG4hH9VG3aSCEEa
dFmKnOxfpijT0gFONnStLZ7YBjKhzPKOR7+22o2zo78vcsaHOLs4EJTjQ3I0gkFK/Jp38c8W/8Gg
+/ODl6S/CrBSrUuT7ug6ipZdoY3hLnSe6Hy0+tE78otXVcQSTh1IKKmZqG3yM0nqAEJE2l0BdP1Q
fancpucEzYGH9ynkbjwdHoU9mGg+DdYzLq5eXnclvG5kz6/4Y8wQFYpFdJEiBbVcUu0kQ4UV1Bi/
cziMPe1N7+rTpSJbLmDhE9t0rU+SIoAVlTgBDBvyu1Z7xhP9GZAlJh+eYlCt5bEWIdSyHfm9lOf+
EA5/g1/HKceb+BRnOzYwtfeB4GzhlSMAuSPILELrtQPtRx1L1znZbes5Dg4gf9AYbcjcxM7FEFWG
s0WFhFllOu/ttZ/kFKtz2mv6fjLmT+O6L6BPLnGBKIM+l4koxHm+LEzrMoNhWecTUZQl7i9zyJUZ
fRykykRNfcUlu3ssLAOS4kzlMnAG8cF1onigFqR5sfPpE7SfTN/MC5C0FdhLnDbCeDWXvmxn5BZz
nDi+zO2lN+HRdnCEcjQAI8nV5ps/dN4ctc5tDliUydSgMK1Ojtc/FpcNpAbkXIgNyANt81vRhe5y
XeXzPbF2Lqbe+elB+L//Ae2VsQ4TYDWneQlsZYSzd98KPr0ZqmNu5w4EQoi5RddEZD7VECHgdOGb
uV5s76a+aHeYArSGeZKo3F6oowVBgGU7gVFnxL6HXHoKaXiOa/8F/jEzmfh7ZSUOqkMAUeliaZcW
vDD5KY3emg0Z0pJuaXM5wrmBn8E+m3jS6v3y71qtDCuhPLKc+ojmWHpifDynLcZJzzZGx34MATFm
p0xbNvBSB086fHuafjM8vQdPrbz8UOA7UrDUHi5i4IYa92Fl8Rq4Lra4C+MUCsLxwOh+MDOTpzEC
SnrgnRXpHefZFtpkHAeuBjh6uZP8eH/fBPvgL3Pt0ulSnrNz3FKS9osVprOVftzaHKIxRfqr+slZ
dxqis1reQP/hZ2A204rfRMjGcIWcPnkTbNQkiXIQiOUrNkEUF55cK1gC0oDtkjOrRi9CJdeAVgV8
ajGKLOZGxKftKesn3ik1MZeGPneKNDmcJEKTnHSFyG+6h9yKmk1muDjFcf228rlWeCJnc4SSL6ek
UXHshWrSnplw/5Fx5+wP+sUbAABdsxZ8N3Kbq/RrM/gTtv/PzMSp60qeXCYT5PHSw96YVGXBWUgB
XB99ACcT7336nDWykNXmllY123QVjH/qnW1qlZUhG065jCoF/nkKgKuxAv0+2JrCBNlfrS0/cEsb
3cYnVzuRInSoqjZBbDuCKGQ8NXZ4pMnIvCBzQ/n2371o9dezeq/hzf+hDoZQ24Dm+GtQ+SY/bimR
I1yQU7sNoqGaDVful6z4XeYUyQMkR1Rer75gMv5i665DYGayhZ7Z57wsessXcL1dXWPWSBzbvut1
l2FkBEIuOcYHMxjSX5U4tjtXEX6NIUaqnGx3XkMBv+y77KDGjjocr0mcWNlkEMLDlHJnHdftPz8D
DICAhpT4SalYtt7hleEkWXictVnlNNCVwKi7IV6saT28a2KSzeg33/visiFgfINzmkSmFQuRCiLF
+IhMs6/dhpyfu7R7AGfatue5nveKKtuGiY+XMQwr548SrIEsii60WttmCdh2PWtlYPubsjaVXtKY
93Hn03BlAV1t3o621H/N44eXL+MXrIgEtuYrImhjgvSiZptjYr9pm5qttdvfe9HO/lhkEdnwbYc5
077ZB/kkk7Xev13piEzCropw3vHJmWenaeE2Qzp+JV1nPELTP10mBa2/m1/yiATD0MJQpQr9eN5Q
Gx0v8iNcyRoOj+Za6G+IyMcIgLnxP1aDEwMqxDZRk+kTMzNEvCA9oCF60WoyFAuklICGg7iUWjxm
4hCbBYfgq2SJh7cSq1ycO4ujP2Fqv9FVyUUhXU0x5fiTQKxb5Z2EBJiVgO2F1NsGjSYtv1YUhP8s
77Iyoeo3kNabvmM6NhK2qtS/QJ7zrbdVu7z3EmoyMpqHnYeoN8AFsKtovmTsMFvp12RmVPB7aNBP
9Vq4foB/gpnUvPF9+OYxZyxm6ZH+HK6AK9fkBNf90u8ZfJc7jvqccHQOcboAJoRR+WDIWzPYJgWQ
q74GyaJmtguS/tbLBFoEG67HnQRkAP4XzEKVVKvY7Z9SSXK01NTAh2AZ/PuIo921L3reZ4eo2Nrs
t8YIWbpUkWs4F6NIt/bVHFTjqNxV0batOl27lQf1bm26hJRD1VwCphiClLT1cqS9bGuqG6lDme34
n3yZZILUikizlN+mkcq22uhZ6SuJh23A4R+TTWoKKMtkn85ACl635S7ktil9uxqb3QoPUfsnJQvq
tup3CtFmYvjdbcJ/nnbXIX/hNYkVlzydPJ4q6Ed/eqoLtqQMi5LOX3o0V9UfRolpM2zegLUa8OkJ
WZS2vujtuJi1MoDf4m38Ci9TXAxZ8doJliW2YC3JOpF51s6ZoVJ5RqeBdtniy6tI9/BM/kvIivcm
F+62nsI8/x8Zl3eyZEAoG4XcuchY6Q/+immeICjmDtBDlqyU4xdbMtfZc6J+yzRNyJKMadvj1A/F
dMQiKp6e4cTh2zT7E0DSvO/+p0N8iAzhhew2fesNRETTH8BVksyLlE2xk1s/z5atfogwMwo1AO8d
1wz9XQI82CImLhIwCEppdUp+HZC0+MbJc1edaPZmLYKRykOE0GY187s3+e1A1r/IOc4gVaIHf7zO
GGpsztkpxSLuloxYyDy77LsCNnS+lwkknUPCkv98TyADZZcgUbshPL/D/1Yjbp7xQ6p36fPGUFEv
92hOWDUBm45f40Bbt2i40ydsOSEUcnyAg/k3lNxCggLsTkABkHomWa6lfWcUlpicqshD83fFBBtm
Is5MnIKqHZO6S8BTdLCvYbnMbc51hR/+StXXrxeISBFehKpkNpXH4Mc4liJmEKXL4gi5MQUklHUY
JzAv/4qXGE79nmdMxF2QhZXOt15vWDQim17JGCuTl+SLFu1wL/xh7umvQyFviTwo5ZmzjwtdTG1x
PDleo0A6uqNVs2gFtiOrlgzpyPnAURfI1+cMvyTduRZDl065Gee3i4XlheT2W9muRhco3VFLNOOR
i0s4UoyAb+rEnWnZdiHd1Ok6Tcl972o5kUI0kUqfFdaS7OnAv3oJ+DKnoJeJQcgLWo30dSRLlnBy
eVlzAJgDNnzzoOC9EvI7JcrmjXNWunvVhk8YVdDXUF26eGMjyIwkzq4ASAuz+De4YlK2jzEbL839
JIw1a3PUsgVlDzBiS5YzAtAEsdUpkOVyo06h68VDRS7zVMSqCWIOvHJUNqlbllK7Z5fuTK6wDTIh
3e5xlL9nDdjF8Cnlsf6C3UfMerQDa4DN0AK3nQ+OXEtKMUVEe75n5lVTxd1xbUb+CNWsW+PH3Eje
WCmWH1xaSfumTJZi++o/iKaDQNYIQv6k3iwXPjpobkknBk42Fx+h9pqIVU0I8SIPjSqdc3iT8UGH
6gtxUoP+Bb62/M2hOt+8G6gYk4luaXOl5E3mEOvwT/R0dDbbOIuRnK/0X/Jg/Dj82TRLZaZzoxJM
KGB07pt2WmhRhI0xD+/KSqIo9zIARCKniYv73ksI5NJU4sUvBaW2Urk/hTF3+c9KtZOf3JB0uzyp
frJKXSUsCjhzWP1ZYKO/C0GU9Fjw5tG8Gyq3jmthkaTC8YZ+Ky8GrP/M2eFQmokC2Ul1Brpm5aoe
r/D7H+eYU8K5tReV6QAzgtGlJXzpEVvo2eeOUtYzjaoEqibpfF2/dypotzeta9XgdvtMI1cRi3es
VQr5Tnxogv7sh2+xnn4iYj94sUGh7t7CUFG2g3+6AmwCfdSros+Ym6GT1qAjEYuc/usRaUzfPEsQ
zO3IhcWHw0pV8EavQbLkMWSQk/FWQTPpVKngvD/0XLiEEC4OXB+SgQn73BQLyWlzZfVpxtdVZGLt
L74sw6i8ToGpGj/36oCHtchiP/Yk9m4iL4Axrc0w1s396uL/ogs5B5KD53UaPdOY79rcx2QDqJsF
/wRvPs7f+XPRlrM6VHNER6awXBGJl3bi2QyIvpLhLVrevOS5KHTxlGALvviEvarmWUiU40Vw15xh
gMon9qK04/L/0TeZNwAwQ43Zz4H1aY9J2V0ryp+AYJI8ixAAn0jTpvaDe+TvFyQ0u2ATEDE6rUXx
VbKV85L9YlpJnRd9t95RCIvXtLXV31RwnxHx/AZcsmqsuKKOjMKTbuOaaLtl6Z1hBApfeM5xdGFg
yMVjM2xf02WKjPYWKPJCZi+MwN+TiuWWb6RA5XJcQy/wXDbi9wKIaRD7peGGjLjTgio3Rg8kaU4u
dxSoHTRyGEvbip79uVriAhDuvkC72V4iNL3SU6Re8EFJx9iFlwEHwhyeZhUpvy4D2boFASnQteNW
ACocA4Zutk2dqotS4RKthWQlVGdG2I1L6954WpYTxracfHHeB60ZH5nSwDumZH26HdUS0CWAfZ3q
OvypJwtLjfFdNzX4G8+VFVKsMcEt+u52OQ3o3hGvq567Ine+fNjDu74R/9BSSJsI1pCzj+aMTy4y
43TM2wbkKpEET2MrD4WjFXHl1IOI4iK+8GKfbjDARuxJACKVdtslvK3XDfhfgjrLToMEN+SH+bhk
UhubITvVfq2kLmu4UTDFM45TOYgNh/FzSYHfwqL7QT5amm+c46Gfo2Ym9YXFwl527nqE6VJfRy4H
keEcP3D0JK3bHfa/UIR+o/RhtOlrvLSKKKQGQPGyLPni/oZ6YqLI0h039T4g+Il4qg4sQE48mFw8
uTPK05BiyX2KNbefwiNtt/U6ln2SiB+XMXZVjC/i6cuUck6hspzBp4rEcow07wAiFFbdbdtHvXJe
DwJ1hDS4cCCuEDVSzo1E30COZljqgPg0TDDoZzBWlX7/9XZzAW2MwjGH04/zmCziPiLOGjAkdoqY
Bz/fFZOIRo7aWNLDbJ5a0mfrJcdehSEWWVGjwMK+AS8OchYF57T4VjthrZzRRj0XQ8bxAdy14DQR
ZRwLMCr9W15bBQBCBv7bfRJtb2Tq67As3beg10sYPH+I6wLIsHK5+S9++B+z8UEkKmGa8RNgJOgk
F6EqLw0IrLYImGaVdLNcB/2/O9kbmjrNuFcwDlLWgXJdt28PcqnGdo8rX06P5aP8lct4cQW2+9QD
yxLaPnvQ89sFWTrt8s+EPgnFvzxIPmmwl8+WAdnp0DvhA3YuBeCbjo2NNeZyl9HqJ0PTMp1oDUa0
IP2CqjDylSAVnYislgCduux/0a9ZxERYLgEW6Y2cauy5oATUf4Q1Ms+WJaI9vY0P/yp7hpQqneXL
hzu7JwwytYLawism/Xfs4h3Jz7+kNt3WU0wgWwWU8upOhcktm/MEjxqztPZmg/Lo5jx/CmqZyF1V
mfhd/NW+XvaLDyEoTQrfgVJD4Ig8wLUkDzu7+9hAhDq2BPmA9aMi3w6aaVZDYVLlX0DdvqZTd0xf
7qwbeVeQ3gTp37CXqHqRKlC950in3Y2mq2x8FIoBp+3wvc6HgIDcVALwIqA0psHs5Lfd/RL++NCN
I6QWjQq938Nx5IkNqzcnzIEHfI4ym4god/O70319ZYZXqQfYo7M8hKw0zspSi9yfo2LU0WVyCrHA
vkgQk8LCexdwVWGoaDxz3vdNF1EUhv4f1kms4otroXZzjM3Vy57Rhz0ABAyhGqzI4GdFtBNPw4Ci
035FlAQTZxLHRtfCgb5k447WVKuLCagAEF45yu9ZEpGX+7xl2qHCI9HksQQ6Q0NGSrVMqLVxlHH3
QJjOQ3EiV7TI6iNsd9vY33Sc/16iAo8chv/hFH8BZE4ir3Ftj6a5A2jySFqb/ELMpHvKRgQEeKhz
RE46uszrG20hyoSie5x+tTf/o0dG46SPX1cRrgrr0aRoWQKd8NPaqrMNUJlz9Kaxa/6URkrXP8DT
Lx6+Ckn1fVtzZeH5LbS06LSRqy78jSyqxI6qjZJmWlR9wupCJA3+HI7DfLJGg+ldJFWg6HQf/jI6
ojehGMueV3tt8/SIExvF6QK1a+0ca1ME0CP8ZBF1bJWUIK2sxrOrLtFgaNGvJPfA7MEHQmon6vIT
5J75X2Vb7w8/8CugSZyD9ThLTbZdhr2i+I5dMNgrLWv5Va/T3cZ0K+vXMiEWN64+bK3LoIBQV7Kz
LZQos4nCMlqmVF1eYk2unN3VA7remXCWndZQRzQtTk6xD4bkYoKuugC930w59NijtYaiDu4bxPgy
Ypr05WMLQc14zpApea1VXrk7TmqSW+PKm9KvDJDLDMERVfjyR8noSC7fF0OV9uSC1/6vlNaP3LdH
l1R6TCwIniXSPVttJJ78ZFofR4j2JxLTN2SJTsors0vzewFLEped1phRFRegHJKgyQfzOtkPu7D5
Uo61cjWDyvXMhyVRS45i1COx/QOcwmyTMPKrQHa61WlA+GdT8M5p/ukGpY+VoWnCJCFrXz7MJhwN
EfJ3Lt2eOG8RtELkmd0Ck2In/q0DSsGG4r/gbf1fuVOJdmAstzWrHtoCCF+g9WxOUlk8KXC3v2fT
ybaDJ9WnacdGDl5nEgzV3yBaY9CgEj+VK/GKVJ7g2YXQ3bpMJqvV3tIi592DAwVgZ1YnhGQXRI49
uus7PzXzmFeo5P/B3SNSSShILxH0TmUBWrHH0JUIW1+IOjg3BPP/xC2IQ9kKB1mk2MsmRT1N/01w
aG/0q+rtdxUGt+5aBkSqv+hfV+Uk52y0mwG702h+71oFpHRISLlpnmgpQ11ueZqCGEAZ1NAmyqP0
YflBLLmOCBrUJmESnu2H546GjoalA8QE2Ue3JAciZgJnwlno0GhAba/btJXs0nsX7llnKPZ9t6zW
i+IpYj1C9T5oi9+BCEQ1eJamYtxPBoMpxRE1a5AJAubQ4vNLfH5LwXegRZk0dUz0tmNWFBooiLWy
vM9HHNz0iOAznTdcY16patKzGbedFPlJWgNiYhlT8L8T9XHXqhRbtsA1WJS4NPKV3XPwkLiUzZC0
wjwd3GcZJ/o00jA6KfPnza1X97al3hwFiPBNa2cuv9gcfL6TcV4qYYTiFpn2Xajo/DosNNjBtijp
wYoB9OdizZmK93PR3IPu2qNpcbX8+ToDcXsCrzrhxLIM9a3e8GOHGBijmwmYYBAaUqhMpl3ERm7k
xbY6SXh28m0O8zmlpitpvEjEZ5Sww6jfre2Hu0bDlb9VF+Fh0eYe58aBg2cXnrHOXE06NMVP/zHY
OTvKgIQOcn2Ho+aYjNHE7Pkg8uwbnSyE91oGOhuuN2xi361lIhz/Uy3WFUg4OvyEEWpX6m2WkBQt
qiH1lu563knyKs3lTchRobJb9CALIVWI/AcJw+aWuPXu3uvBpjzEx4sWLHVVnm8Qve25oNhBOxZ/
48RG/0qp8NkJ4skHdVg2HcCqYQW6VyEpxVyF7o+vkShrWQ0WulzZ2H6SO5ZBo7HsqBteDAPIig2J
ZH/yzzesrtR6PCM9U8XX4tBVanW6xMKBhSTJqLLc5khoQztZq23wiUPCZdzEFQKGyZkGlrivAzUw
9bLuNvnPYydQ3AkfDktIpE4mqY9xvVHbZ3adwp+tOI3hO0XSQDNhSe20U1vkn9VWxLbhryd4sDH3
/yYIm9Dm4c3Qs08NhyKM67gP9R90H6Dfk2bVwPkcZOO9khds4spwsIgiGUjyNOX5TLTAQlBzgqts
zrNbE5f8EDF+FRrw285PFFCj5HiWaLFOpbctly5flsNrht7mOacpJl6WE6DoTvI6Ny0NPVOVNuoj
smSXb8GFiujFROjhjaHeSEQAwJh2f9GBTL0kbgJZ6QEqPE1/CUetLbYXOA/3FlZe+GCKoV4LWfNw
qqgVHYJW3A6xr8F0kcDZMCj/LvTssMBBJbFy53yXksTEKvhgZGvdAFODqRwWB/Z3qAnW0XngL6dQ
i/p4kar6GNZPJ2QgX2PWg6rbTgusjE912K4l51pC9LA6NMtL3mFsc4Hmn7Asm8fEUSx2FGyAiq8K
DoNN2nIf1vZTf5rf08pjBxD4T5RqZJYYyYIZJkWFYSVyCL68LOSf514P9zqHIuYpRjAc6tPceXjf
iKU4LrQaIxk+dWr+9ITK7y97/kVDg5GNjCC43f0VUXfMNkO6BqWDnOBr7sBsrjemjHTGImo4Dpkz
UQxdBZqQsb8hhyziPekqSBsg7lKv36O1XumxYdfZZHLOuPcAMPswNqv5USXN/JDzg8rmZXXN80xZ
7Z3+Hj91rMIoTgmdHIxfi81WLZ4h0LrPmHce0eto3bGGGgDxmDK/JnJnkXaBI2LJiEjIkWIrXftf
xzqvSyVJ7bnXYjZAU/M97xMD63AeIIF9BQmfkxg9fNU9Mf1+1MNkGW6XJB1hucG3VVYKMAKJjzmz
3r442KPJMT/wUI9ayGnIh6S735XT7lXZLdTRH3DHXxo/p8SBiBI9MnK1kkxp/S3SQCpAHti7M2IB
I9Myd9CwP3RhrisVk21//curV/kOavNg25HkKon+6ji4zCEcQykhQRcWnRqmOOZaKT1Z+/edn24M
Wy/WHCVA2yXzDlmL3byRT5kpqFp+srXhKiZKb1OWTChvghQ80y2k/vTHW/gBJhuOKG1DAAzy44lJ
lAU1oxHWa/nPiqPZ4MP6mjNL81RSF37Dprm639fKPtk3vLgE8c/7ACYMysS38Fzrflo03cHYbWgG
q+q+ee2KPovD5by4sA8aVdBPUoc7bOZXXs5nPULZ+Dhhpg07+IWN2MkiiWpyHawNI/50V71PZZ1b
Rzv7NTY/sBOdvyynVhd11i9HsUYGq0aKH/f6M9FM+7WtTAlXmJTmzLF/JXmkjXdcYpAEYC3Y6BGQ
3D1Acy3BcsaI/8X5TmEhxM5KIpWxH3noL0uL4+j+BX7l8ZvzeOdoxkCvSkCDq1mh1CqQ6wfewIwO
B+WPYJZE9ijNANVBYhQJBKYULeOJuvtrbou0sHkOlp2DV9VK2aUHi9vUp4pD2Jt6vz+6RbMDm4tC
PNt0b18Gu0kjMG1KlJpjGUqrvlopr7MwibGLkB+QT/wYHx4q7fYQeeJfATlZsvJIRIB5LO7ZbWeJ
xRBg7ghu3IJTPFAdePBchhIS4wyFZ172+U59SWbP973uWvOA68YGyhQ4b/5QQNaDTBc5dd4aKH1F
AJhhtRISwJV8cN+vLSE56esqjraplrxPM/gmZwIW7rHDnejDdQlKxxiv+s66ScKw75RGxEgZ1EaT
3J08WLujHdajX/MUKeR130pDC5u5QTDauEdZ8j4EKrp8DkZ/FEdCv2MSipgmoiHOE4ZgDSpdjXlY
vD2RAN0YwZK4Ay8jvHmuL9O6OK8QLKYVO9xjhSPujJDnHaXL6inYQ1AzRgmkd2e85CWOAli2tr63
Uybg+wxLmiVeWoPHbq4xZUao02z1KgCN4f3uab0WP67c5VXLMIyqwR/RXsF9z9mHLUrORsiidat7
FKEQYLZ3m0qAE+Xw9FU0beenXJDxCeDjXQ0z/Hv/odU297ZI6RCGu5Tq4RUQUc1vcLbQjR0MvmMt
HbR1NIPNTF88MPeUIN4G+B4MblmJoGoJZx7XOViEXXF6FHgYe02QTNo3TPWa89Scfh+yffx/ALnc
V0OX6VPzAhErxrlpSRxRAycbaDfUajF1t60s80pkGsqYinKTT4+5ZKBff3KDTrPzduhMIi5DlA8i
sWxQzH0NqeQFNfBJywZDcTHJ7a8EwtxvWe6YYD6ndVy3gbmM4lGq+zEuVG0pHrvdUex8ggvUW/82
akM/E+vv7lZRK2C8JLqvfKSnG0CQd5Jb7/xnmf1CJvR786Ll4iIe5maTW3yrmbtmIQDnO6GoGws+
cHSGbA9NaZJWke4F4zAqINc+ge6ftBtDO5SVMoZh+wB6jRe3F9Ve/dfjROE/WE+fB7dJCnvrWo+a
x/4O5ezgTejY6mNktO3NdWBYiz9ljIO8WsZcPYME7r8JELMX124pyJimxrH2gPh7KLxc680PTltD
YOv1UXS5RAxUe7aKkJl9y2Do+SLEsYx+W9qjVa+pMP4Ly64kVZIz8EEKeTyfEB1jOdqxFWD5Ypbx
WWD+MivDBk8MtjLXRTNeGUl7NhmODCJuWKAJq7sTN8APYpUYTmBj4sIi5AnfdFiDajJjbGLWHyCA
MbJi3fGv3JX1hNBlWTdTr/U8XkJvOSJmyMiYoPzNp5o/I861MVuxuEZ1Hk39+pgS+/TdklAMmM31
J/iAxR+19MaAYmHUN0tqw4Liag/Wd2ZIdFJa3xIQqevxDlCa/vmxX75c91rYvoiq+Eufp9TyGQAJ
osTgWk2cvJIJQ02KgonrGqXj8pHYvHwcfKpa4dCY/LV/gsBfqBjxfGE3mZ61G2cSsJSnB9wf1PzM
/bVFEfwYYi683+LNuk0cuzXjuYqMWClvmgiN4LuVBQhEOD0VogD5/Em2Yg30+7f/moS0qryvvrMu
NokpvUzc4k8OnITCdgq7F2eJhWGabrLx1T59kfZ4E40+wgy27fIkBzJIhpJTDtovl/jo6ng61cYJ
wwkDm5Gk+XLVDX3L0BoKiEGxs9b0jDL7fFzwimXDAVnLmyrl7SemVBlMAkxVMbr0HSkpps1useLF
YqBiE20S/mYhYWTJnMyx+DpZJsbqBzbXTPfKqqkzL3pgJXdp6bkb/qacvhaxK8403arjQBshOWgB
jTU/boy5Ly2cGmJuulcvjTJWe+BgmpG4y3TUZBHe7gB8ID+tDkMJAMZT+qKoywkrEI+xvCPo8QOJ
n1t6iUBQqLuj8rBmHiDNUTiHVZLU0EDu/Xow5ISSoQtWnVELIVehJ9HGs8eVrcO+A/rUSkMTE5Yc
9oH7TMBVoO7WFZXCPwSiS2um+YVtpxQP97IaiD4lpP9Jx0KPUz6zFArNHPW6XWJgpOO/ucCUsriI
Znn9xI5SbU7nd0N40IBtbl2GgW7SYqYukCzBPJ1zPTVDvFInIaJbjyWPGMLXuRbgxea4KoMUuHMp
zQzpqeR9BqhidOx4auB6231iIyT7uFhQOzXe0V9oXWYz5dK7cb5USDUlvnGF8Iz5Xn5deH5AelAd
G3LEaJII78bLxOjZiNeja4S6L2Eyhq2+nOsXHuTJoCmPXYNJtiHYBLecEQUpH/5s+Hz80ZoPqZ81
Ibz+C6Y4f7+ueuejwqpAxqV5tbKocMku3R4rhYxQz1WfCPz4SXjub+qMT4FdENTHLcuPiJA0+O4l
jrQF+K31a6qtAANxhIqlF6HFQ6hjIvU3EY05NTTirdrl4SNa+xplXzeFakiUrfHRXC6STPlDWjkk
tnL0uAL7o+nFnw+nXL/27wyEXv2wdHvlUM7S3hmJSr9GhvqW6lEs5JsVZrA5H49EpZAIjipq+F/U
knV0wpcPFS5eTu+6Er9RUvwzrWOBTBZjSQF5D1yaefCKIvqEUno2L6CA4Vciqpuc2fQI4/ulUMGh
CEhUddocK4S9Hb3vIh9m9TADcK3TlARt0i5YRgKmEXJ0b1o+RwDSG3e0GV+D4tUzbduIEnSHdiCv
anOhoP80nNXtYwqpFuIqKvwpgoMJ7irKugL0Q1jwWxoxLJJAqiF0SrqLepYKpRa8FZG1orkNVRCA
tvrW7It20eNFW9xtVcca27xNRYqdFhyEu/uInDEueJbkXCjnPhB/q4x593YXQE9Gvsi0F9IjHotO
CvCX9c9CckvK0UI3qKm+xZPKqYvzHyrSJ/JTRmWH+RgL6HB9l0jhdOUaiTMxVnOzPPHnfTc9oBOj
ZiCiVvEMIwAge+ZdmOfGBMoxsGgD+hmd/gTolxuw0pVN9yKfvG0zpVn0VysU4UBrvhI/T0VaVCPc
F6VYvUgBvYDAUHzjumCRr23Rt3HPLBZ1L+DXeD0MvccXFxFxosB1A+Y4UTygWbOqOwhWPzSG4Kh2
9s31RgUDfXMgW6sE6OrRECtc/ijyii/XetS4eWAT3NQj83y4kNBILs9dwCMP/4HCrIT858d4rx3z
rrkLgT0cQhyVxpVA3ZX+dnNHhWym+69KOJ7f0n1C9Pcv4nI8N0H/2/RcEc3dPvPXoq/LCChOO1v4
UoAAFE8IQl0COzj86ExyJIe8+nlRyWeT2j9m41VJ6bz43Y8uA7b3YWW2+NHmJKR8LEExNSzSs3UV
RdkUGEAchJcEQ9Ea7dxO7XHWq0QZppXxT65giQebPw5iKD2WxcPTeDNyaZgDvAxk2DCOEmeNa7kf
l9/qWnYGyM5gaPrEULO2Mfof/I4/rpwP/ISE1nwVF3gAqWFWPo+LyjlaYJ/uznWlPoZQ3sDeMMDa
WJUHfBxQZcQMDmR248G5MhB7zR5EUWTOHI4DV8lAfRZokZWRmLwB2LrCqpev2SDpRdf5p/c+2NKD
uLCG9Q2Tk+mQIBvUQubHt5kWNcMWcKhzN4ORmymfPmYEIPIfhbKoB+z31iolQvGTTDg3XDfYUJD2
ahLdpCPA5t9YuHJxPmHgQa4lfHlWThc7wHEBB09o4NTJYBuNGGGFA+9iF8D0VsnutJ5ncBcQEBkX
rEjSQ5/j+BZ5xSxW3uIQQ17OL+CTo8FtWGzTa7SIkmWI/D6mlBMUEbspeZ9BRvAPcuabGl6Uptxz
P80/9lA7cvTCDwTm83ANnbNmZU+YeIHl313qiOjef9dOmBAoFWGCi3CRLwGOFjJA95zwEsGgczcK
11hvQbcVQ0a7R0/Z+3SoUwj98dKLRYTISoVfOdKnift+siJ825se3XonGgSJgyGRupXrYZOsZYsB
UtvZzsUYKp20a2fzTmdnX63eulfYJZltPSAC1rqKRLd3z8IHM9lZIH/2U3mWLrF2hHa1/UX82ZQP
9etSKP6h2S09Y7huDBrUzq9RVlEDwquup16NZTjkFgNXVwDH/vbK8nEnvZEvYFr4sopn0lTg0SeK
WjRPJEm5oCfYttikOpVpMR4dQaDGjRuR5bfkB/WAwQP5TUxhJI9M09eejKZaE4p1CvGNwMZi9bm5
ULX9W32fTlvU9lLcoxzAEHrTKQSeVCipVfviUYp8OyOIeu0RCU3ApPh6AbeMaKNgZ52Is+8Y1cp5
1o6PBLHe/1mUGjpLkMDYEHcxIxNGVLMrTo+PwxrDBzndnFc5Ln/Kgd88s99XNl932c3I/LfBuNpE
UDJ4v6DnQGF9jLF0y0fzQ2yGxL9XAXpIzsHxxr2Q0GfwPMSPMMknLrVfavioFZZmgjnlIC1AEZmH
e3Ntd8b0Ad3MbkgFH3g7SfPW0Xi9zcqWxD4JO4XzxgtjDrfgmwkjv4poeEh4e8mqYSTqnkyY2oJN
tkVJUdGPNTu810YqVVkoPBpTOLVv7wNecUjFvzf2sD5w7fhrhw/U98g4cT99w+/TfsxWq0W/26xE
s0jOpW4NH/wWcpRm0Xh/csV1Npl5UcURBMCQEooZGK0pkQH2jylSohM8/7mQ/krkQNu0Gf1TTFWz
CifJpHvLc6gla+2pinNYUCAR4nvMzEUSao3O2bfCT9TVn6hN2HYPWWVOjtEndd/n9DaKu3l2g/l3
/JbkRlTKHmv04KvKB8HktJQ9TskkZVucVgHjZGDxte7QmUOXmHX/lS7wCErnUuwbIb+3FIDYKpsF
EjJ9rQO6AIoqQhLwLqEPr2Dc9+weQrzbzCp9W3TMF0oNe98UJyRDuAv3T+5LCDgw63QKdKeW53c/
6ai99/yzcEduje/wgFcdm5GZl7sc8lb7b/Rxh2XJCbBbsyaW5I4ndLfwlnrKMV02pMPpaXIJY9Oj
pj6m518KWxeehpzjEssGMvB9Rk/13QufoFUYVrF7tmHeoP7MpY77Q9i2CYl0YZI3XFxo5dtC25oe
dfL5/TU+wqxvc+3w0V91OG+/zUdFciWzpZxVAXSPJgDBAEaXIMCDv3pr80QmO0gXEGGXzT+EgidI
MsyCwFP8xvTcqD+wkgs++BIf7HwznOuyNxY79UgjUn1uzICVvWN9TrHidD+4PKLnGcZK0Omd2xRW
DTnCdEN7qKOKkNf1xxCEdbQ5inODQQn93Kb9cfxmSav5iv0JAkVeG2Ub7Hg7GGrOPerbUjaGoaFU
7nyu/fEebnt0mFpYwL/KGTg5KLz90zVcUllHzrRk3J0AOrQdKx59eagcqBno8zMkkouhhzNZKIrP
Hs70kc6yP+9zxnxwgu3BcJbCJuH6XRFqGxUoZ2+q06uZH1/qpJExfi7kz+9h7HOdX8PAHZPk17Pz
6Hd6XXtkzjSa/A1gh3HbVp0bHXmVnLjC9Uw+v2JUCQH57Jp5qWMIVFkA+5D0w6c1d+z0VFn7QXdN
qn910JDpX5uParSp0Le2nFD0gNGg9r0UYZjDm5Zr4HO7cHA7qMt92KWviFOuhtqOgQk3LNtLRvYp
ka0zLMOMk1cff4yMjTLhyhjGpkLT4LCt4zIEr/EFG7R1rRSL5J71jcnpcGxi4Yw4NUzTPYu6xuQR
q3sUHj6E4uH8BLJu971H8oL06D/UlzP5Sgs5CF6V9tS920tN+SPWNYTa9yfBeP8N8zMuOygDxG4X
0VGpGnp8ASlZALzJnzG/knKgqlpc0bDeoPwGtmh+6PJTpM68Tltj5iyMvQKrrKnHJFPDEyAk+lB0
lY4Oyk+LkwpSSSgJJ1h+a8Nbye6hNmxtGjrhNuZ6Dc8dtSjXJpvhfdZeRTx8cFUcvLciJkgdmj3C
gQIWG6JWukRlth0pCUtouljojcRnOxGgRSlfXSUVXtGhja+eqgleEsgEX2tiRdZRlTZDyzG+weEv
GDpR570yE8TnjHBbyeZZS4ghLLFClp6HXlTXUm0lcvI+0k4NuXPNaokFb6MTApouNwd2B6QxFMvF
r7lCJcicMaehpwKg7oCL0nO+UI+84Wf7ODVkkpBgn5xzQ1CiSS9cK+r3/M1vw9FBdB0HDqzVVEF/
hjT6zlG6SUSHhlDPYn80aivr7Y2NfAfCfqgrhkV+qdpuj8VEUEO/pri0eyFcWwju5tD4GZl3Fx1z
IJwxWAnoULnLx8iiDEoi6dp7j0T3llJl7ELx054QBY0wP8+PP2j6UETmDSAiyAeXO3RXW0/8eH7m
SudEr5LUr7DKPWYI7h5f3bc5ggjP2DkqejqIqpbjfx+BEz3oYk9PI7OkvxF7XAXgZrMo7dZuw/3e
ZDUBcx+cRG4xTiGPv9DZ8xsuavD6y4FqM6OKvLL6cND+ocUVOJkcabPI1KLEll9RjdcBsDdtq4Mk
2yQGFGZ0fvK+w0IbAAdZUZOEMsaEdkfIY7avrPG6/gTvm1BhKqHPl/R8lYasM8BAHylOjJdJXejG
wCWYtsmJRnfKC/QUVyNKx3sNzbQ0wjKQUnGNwp3qj2rWHjmHrrFYSCqHuVcC2OT1LYBV0e+gqhTc
qToBpnRPxNcvhAcGjNkL/msFX+Ai8a+j0NIcloC7eqs9MgavymNtFTj1zLCQJfKcoUmLkEz1pvf8
eDZTynRMq1VXlsR/xKRU4W1VoRXfguguYiQOIrnPQNExrw7Ih+99jaDGGenwV8WpoRh67iUZ5gcA
kGVmrZ0nKWa55KDYPbvS7dlA7JH62X5/v8fqXQMLFzoOUyBwKyrZWbuhZj+tf1taHwHtxrgZb3d0
AbeeCPzoJDp3sJ71URwGKcAFMncufIZfDyRxcKqADv2c5HDrUQ35YnUZSNq0F3T5lUBk91Fl2D0m
1OsRY4AYVP8xN8mC/kGEELF8Ym2ya6/IdWy5HAhjqyZohkU9pXS1fFmTM7Fp5SpXGIiPEV2tvvAe
j2ZTET7KZGxrIEBSG+WdHNlucPggHk9MF7d7xvTAEDNCPM9JgjqPJJ+2PO4emBHGQPKzPhOrvJmJ
VU/UE+6YYx2J/aa41c0jY4q/phNeyJs8BxnSgDfuqPXlPrztHEqnbVTnmJxk4Iw2fuzlRdBap3og
9S0W5J1bEpmt1Q69KJBPj0qRadJZKwTFghPLrILZ0sLF+O9cXHWi0O7AUt8QjuDHyvzI0R2t2SLR
2NBnRIJJmXv1dnoiUHUJ01ttaostLdYiwUlTbJBXcHa8icd3Y2X7iHWKCImeLcbIsLKWAl5nqNGT
YJ1UJ3LJoC407NGryH1MnQfzWxUum3utEzJRwPfL4q9aIutnoyvCgxz0mL3fRKcanSHMDvGTgAqL
SJowMVBuyXoy5AKr8OkcwGbFO8a4Do/9rmfFzqg3Ub3jesdb0f0pEb/VhIxH1PGwYuUoQEx8medR
EHYZkoXGN8GFpLkBqymaqo/nUe5W75Kn4Dk8z34Nibxl/lqdyqHQXZhoFbeWBsDEkpCdgKUhcrlK
LVHPJH5ygnkaTVMkUofhQsDyq+sBZjth2wJG4rfosN9+1r5Zc27JiDRJE5+cj/BGZCmRuDe4N5B0
D4ba6RTinB4NxvZqZjOB48gMqyVAlEDGwtaCjHkbya4Inf+UGZ8cEPjk38wUC3tCBNOxEHmQAVAP
4NsSals43+5UhiKctzzaB0h9gLXxarcm2rfdPWbpX04zeQMCvNYGCE28ZKtKRrRoeIfAxtfbwmTt
pzZ7T9a/ankNFewMT4XoLelxlf6RbnvDCC0eiamKF3U2nVmrrhFUUr9tgDIlzcBMzOopDRYEQW5D
jA8pX0fYaDUvnInwIToW+u7p+DmjNTtHWEd3EwZkRNDTupJx1FgGMQ7HOWxzARdpoWFmO8YO9ua0
bJEA8N542/eYup0r4p/HSAlOVeCbSLnpDORvkiN37DcS4cWmDySVUoZM8Ru1Ip60NfqoOx0QtUw8
9Cp5zLHmnZrPlfCL9a/qncsXLV2WbTD4XQpYRlUKnmaEhY2qxG/m+NugaPiTTUzO3ScwbG2IJ5QC
zpQv3wf9ypeJNccLc6VfOb8qqDVau9JQRv5+W4HFtdkZSicidPAaPsjz0Y+uoKVdp8hos2AInulq
E5CyZiBRlv9CsN1CRRhvxWmuqmUXEyVqGY/LUewGmI0TT7rFrC5zS+5o/3gZbox/UAh83M59oPvH
lvOt5nFEOahbQ853uam3W+XvehiZcN+0yzd3N9X2by4DV+cDnfKgY/CsDyvqmidoF7OgxcCeWL5n
nVEyPHtAh5DJ4wlfeeI5kayY67EN+Fjru2+z8S4nY6MeFw9IbyYIkaRpMbdu4Rkr9UMu8q3ms6d7
LarpNo4egWtFL/Fp8PG8nd+oWsIee4rjpj5zqJTeVK5Z5KEsRBdD5ZGzybG99feRmqLeYi32wpnX
VraZ5i2Dadd+CA1+hKRXpD/PgbxOQ6ihWhOaUzTMeJ2Mnw2xlpKU4i2A99nrtn2TZeyerdGNRfR+
P6GF7s4opFAAIUN/znQIeXv5o4vRyM4Qgy+wrXFE4JBNqqwb7ifSA0s6sHtSaD9TaPp3GluqHMcv
l2CQNs9FiTgJvQyl93TUjd9eS7dQqTFdyrz2Y27YDz5GnDcJnyauJI4yyu93P4p28g6n5vz4NPP/
pVIMa5lw76u0UTlUumuma7Dg5qiEMbF4D0INWGoUEQyp9X+iAtWngIpvLsjYVWbgFEMmCwrpc7Tf
brIYmdsMT4KbWXu07JEchGGJuWAlx1sztbwveJ9r8WiAGVLHrd/vLl3A3dDITenGHqkWlmIr/jZY
VH+uzoHvUZpRylBewrd/H3sgJ9CMCmU+i7ZpjPNaA15KdEtO+4ON5Pd+WHStl0SAVRcZUAMH+Zs/
XYFoiIRp+nmgV9ZJsLRx517RZeM3lcmRpHLdBPODNK9nti1R88XAWscPWmJMKdOFgjQIjNRf5XfC
e8Y0XJG2jpVXYNJ7NPX7IDKw9fC37jHm3b93ojl1Q6wV8ZuN+xuTyGta43+vpUNr0eWVgq5JYtEO
04b7vLrFABsfBXd/0y/YsgduCQzWC2DGu8k8kVheIVS1f/DXBL+NHJcXosDMcZOZ2EVp3IOEzQB5
ANn7/U5UTR92AhVH6ZURJjJfwFECBitS2u+rk6HR+4e8hOcYGjL6lQcJOX98CKpI10UKVwOHVZVA
FDVxusy2I75HUucKGpAMu7PjRxfww5Qw5x9ThO1fajrh3ur3aRQI9J4QtXVVfyIiFBULVPdZlSN2
H9y1BlsZ0OGwhuXvhcgL01TCs5EJFrYB+CW/mdhzqcYC6pYT4o2ux5iIy2UD46fFAPBJzy4crj12
oBfpXYukuypAy05XQK+xZN6CPDmPx+v7+oXHfDbpooW/xRpLpwNDHDPGtkg/PyvBi9w8kK5WSYmj
L+W67HABvynAZTxAkvauG6FDckryjUhr2bShaBJDulyvpkA2q34Rpwu7SYgSTKJzbApoGlubiNtA
lhxyTTWn6AZ3ShLfAeiOPkzbDR2Uex5Il8EYzSHva5LKv3GUX3sYOAaFgrhiRoUXG4IbLIrqiplb
mzHbN0a+kcKQd3EWMUXwZupTkZetPZUrmEMUhCMpgZPpTh+KJc1kp4pGd/e4vTGLiW+Uxt5Mhsu7
aKWCxstyREJRiWIEt33fTHM3xc04LU04awtXdJgF/qLZrLt2SMqSKXkIte2Ds2QwzDI3M0vKjm99
mlM+2BpyzyDkeVox5/tD5Q3RV3l+kmO/f6WXXhMHBygBJAjx572OFbQvGF8yToC/HCjZezNvk9JC
+TClwt+cW1j0Y+axJdgNnxZHV1wB1rwZrbHIDZS9fSP4bWhSw96R7AKESst/Sr1R2OfhbJa3V7x0
zHm0HN8xA9z9lN5djorULpF448/Hdwp5ApfWG1Vmbemlx6rK9OU9VdPFB3t6NtQA5QQewF/r8LqA
NAhQ8KzQKpu4nTYdpkFSLhpx7w4bYm+s+Kx25oTkh7susbEV/ryvXCvNqL1tczId8EzlOnICGcz5
z6QrOAdu++jMcviS62yl3Lrnq4EXsLVCTY9Cj0sp5/Ane/rpbm+GCz78XqBjOUFnIqo1sVKZpi3I
MbUI2Nllh6a0fdBQx9eK9v6nAWzV+17SMCruezYfqdkD3QfcTAGfZkR2z1fU2kqyHmKPOM2nbwLh
AwKJvzqbcZ9muNy0cDdhduXVAOH4axR/t0u/21jrIsCqdR4GklP+orjeK5N/DkBwk0nqlnNo1I9K
gnxYPw6/N27jTo/nq6HQU41r0phpJH+sebFyiOaDw1VdCK3UXk6w/y2d5yS/fCIcYPSzOjCYm4B8
9t0yw8JR1RaquEiPpZt1vBNX1eR9U84oLBX5NzIAi5voPAjn3v2WKVkITlrCwuqfkmsm4UYNOCTC
v6OtA9WDpztEj3hn1PtHsfd1Dh/zeuUlniQeAJgYfugb9/TiX4zrXFuPr7AY7aGIFSYWcVJzdkiQ
gsu6tlfElwCKAA6x4YJOhkWBiTknRvPbjVpygcDUSvNghsqoec2Y5BfwNY0ZToYEtKzjiV9LcS2a
+GtiUMbGIdgayH6bYNvgWgNBxX4MKXvNgMxnqM1Noo/FlvdtO5WAHggFl5EDnUIh7zD1VUG5xPMP
z6g7b7uc4EN2+JacBMLPfbFpgnxQn5/XQ0I19pwceJ+p8NAyRNOfK+hgS2cyrQsGS4Qx9Kaf66KZ
VyviIluoSY+TofhpqNJ9CAxLt8FHyQq0K7n1zeTP9buQ1LyTfSdI0bf3kGRRICDIICc1Tho43UhH
3Yy6xOikA1/y2UDb+nJniuE06vsdxcisKPr6DxILlLxWLm6j5Z7POuCrkJB2LTH29ixMKuUQWic9
XSDmI/2xWsmy1EsS/JLJmtdxrBJAoieFIYgR7uxFW7ZqN9aYq8QxMBMASPtjjoLydcgvW+yB6Lxg
OgzYyP54SYK4ZdVOlElENaLdJEudoWWSY0kuWyRRN6/kiAxt3gNIGzj96pJJs/CiHaGZZ8USVTEy
H+3n11TKpTSkRcbqAieXcuy58whiAMnGbc0NlrEmAt85OpJ53HeLdXtQ66m0yNxFgvnhlPNVDhXh
6va24leSIWiP1RUZi+rrFwDkFfjOizxNtVtTsRsusHAVUm4OSs5ZqRpi8vTDotojUWfzhgaRCv9t
cYI5MZqQX7kTcp1nKX8BtWAHrY73hX8dr4VmBn+88rUNt/NSrkdOJFu1V5Xykfw0DgX6xfOUCguU
WrrvtwdL+RxGbk/uXgFUgAq0S7+GN2gFWwXjaoNTOAOwgZY6uFpoH2qEtRBPe70O64tmzRvIDZv0
FpffPO0e1e3k93OVf0iF5/MtHiINFMJAN3k81albawK1Qnq0eozalUz92OXGu4V5JezonjGxkkDj
SkkM3AKbBHW10snbFqbN03OdfSkG9rWJp4oBlSSU2O4OHqwDEdnvcmZlKjcbA00T8u7AYtxHMMF1
8GwUDcNTjD54o8F1oCMlIEfuf8/N56/wnnMzNl8fvzHAgsP3MavJDzTVfF3aIBIDfvLEQwMu2gUs
mpeAW/ykD1JaOGWaANS3iXkY3E+ga2Qf1pfH+aUyvY1CH/BkiTp2aBab+H8qDCKLobI97anKktKk
IauAMLX9ERIKHW9HFkvWySLkYidzXJHGBK9xtQddiNacrl3mXLxnt/Hd8VwAtpiPh3ck9oqZaNyo
W3bZWPIkQH2YWO7qPQzQDE3YhftqQ27bA+brpsLMhIto1aVQQtODhN9ayJqZM9BeHLNvK1uTYK87
3OgbFw7eu+qJIvnSC94lKIWoENEYPktvmiOqn/zdQXZSt/R5CYV4Z95lNhd1rQ8HLwFeuvZwN8rE
YiISy2yfMbqjSTzuoYmdnNfKiSM5GMmRQsJQl6FiLXcAS1gvuCehZTN6DE7M+GTfrxpUW//AoX9O
6dIPozBH18hwNPQkqms0Goa7Y6igdCdQoIwdjlmMbOOJre7Q8QxomsUancLUr7KAvcmoazHV/cbz
Dtq5JoP+jDE4/brXK3wBwXW6vIwH3nxNNrEUZopu9PJA7ZPLHTsRU0N6w66OQN+EH1PckTyyWRVH
Y/nayZdpvb5rGv6bWdtxlmgvBJWCAedQvtJhdIweyGZzt/beI/88Nhx1OhTEszV046zvAMMzDSxE
Eh8+sb1qtnOXbzhv2fXK58m2emW0AtMdEcypz+TifNavErGc0UmV8SZcvq50Ia7xqSGDOsxOKCXL
iIS096KTAzZ1AIb9qnVJFVq9HV8jfBvMsJI4x/Pj1B6703YhE/M3IK70xMfvlgAqFGFk5bsBtkGS
FrrLRFXRMFszrGkfC/ATFjjvG11/qjvCHSuCY7U5/VKMUN2w1Wj/Xc7ikEp3h+DD59W8sbBUZruY
ndcbyeiQXv6eyfGkW/j+sJPbirTyi+qgF3hmd80ledEHJtI/ZS8dQws0OPCcSxQBElzepx4IJJNB
FIQT0J/ieFHM+ozgDwCfnIpum5nWnrPErJXilHlyCHO/rvdesxrFThBPwtduc/Q2YzZAhap6Fg5z
V4VQrrOXVNdmTa2WwTpa6JQB1X9FLhLHBPYg96UKXqU8ygjXG21/AY+5WmcPiHXA6pbPvNTMq63+
Vtjb+vraXk1h4X1Qx5Yod2uJRBhMgfCGA/2h6rAJfak6hvZFTarllnU3qPrOHg4twTMAocOJfcuj
cm+/PwM7P5U+m6Ju+tfVST3yasXBqgQOLxbxSHOM2mzwQs1pG4xPN/1fp4MwgPZs0PMz42oHQlL0
kQ+7GtgteiJzX0cys4ymY5irW9fj8N4fG5T9YMopmfESllqmHT8a90zOLFLVhta5Qhy5wnCjH6HP
UEpyhcL3S/EVqsHuUo3XumdVlTXjQqRraYtlFOWfv0VDer2qtZ8BXItexpHmxuK3FT/4qYJqH2hL
5LKBnkYkrbok2S05v2Hy51ixvbMpusz7wehCafIDLujUdBAe0/xU2JsgdYkCQ0WyaXBqbSEnePKl
Tth1QxfT4eD7+1q6Qpb+X+Vx8dpLYFK5JpupmXDR2nlqDHuFrAvIuMCochVDLdOuQzsaONUzFJFH
Drw118p2wyIR+w2rhe3NKYFnzBBXCZEro40H39delQtHcePZ6eU+7luWcsmQqbNnHoHiOEgGrcc6
1BhpCFIIoXpYauX24aIa84fjLpyW848Y2xb1Uvlsgo0k2I612JqRrPhCKGZ2X6jkh8S1e4gX8Nao
HIPxr4mFQOX5tCTwnuGslV+zXUt9F3bNqZZSMe3UG+DEjemFHKyu/dfi8sHDVgVwymeJeCsWQeVF
qgakIITGELcOB+Ow02AMY1MbEuVPuaofw8dHoyqfWRNfeTYPlR0WDzdMDj4Pta6gnnPSbpzhS+TX
it9Mv9qagJOujYZq7X5FsYw3Mw17pvg7gv4vZ0hxiYix8O3shxxXggKcwYZ3OHfIBS1NxAwX7jSx
d3KZ0TJWNZ4JDrb0FpkpnOIjm074fM2QvAjIu9+SV8UJJNl5cHfUH+TzU2IHebe89xsd1m8tNbqd
px+XcZgr5yT/HVy4VITwZzFWaell7nIs4MLXQVdhATf0P/aaRhSrNxp471SnTJwq90hNs6RSUc+A
t3ps9xIlj7Ut9Z7GuI2pN/Jz/R4vLF7cFXUYWXqWZl6jVcvAKxuzfelnxChukalmDU9+2tpLnEI9
kilTL7J9ciCCveUkBCU+IGSfGsc0IOzB7Anqrga+yEPwCQWtPLZFvxnJj6ej5otmSwOy4MEv9H20
/MYUyxuvWIQHrJOS2rvKhvdKwmSRturzIt049DVDu/xo5es1lejhkU+JHqKf2l6Q+Kv+lsYF0INH
NJamM0Vw2ljik1n53Ao3S37HlYI3PA1Vm5O4fghAT4gmED2V3eCfI4oGzCTcIpDtqKhwEs3qnseS
F/xFdAEoiyvvzpJ7dGMCU2h3MP0AKaiCLN8PEbhkdpiWqe7Up59jZSMR2y5T7xEdz9LbVAyopPME
SZDtw0OGLf/yRLURtUIk5/Eu6O/x754Xb/tL7i0i9mkGnikHpwp9XVfjjJ51KE0rdaOw+sDe4OI9
5u//bFadBHcKqFFI5gr/1d6nLhFryTVZO6158lOtmdTDBXVNOuM5EApni+6hhWnNzBPRY0i5uHBt
7z27qkUBVUDM8C+Jyv1AJh7Qjio4cETlJWFIMOq1OATsC76UmdYCu0oxIaNf6bWSg1Mx8mAn0odW
aUaBHYXczq9v8mu3F/xL4JO8DCPwbWCEJjqZRReLPUFPzoMIM5Y1nz/2w7NnG9Lm+GqMQdVrsXXH
LSqb8FkrMaEH5wPB4KjfJnf5a+KPgMwqC4j7CPiWE6UPBwduvTKkXyjd7rHz0AXmvsHymkjEk/9G
kurOPTkPmQtAvxGOPn8K6DdiuHgRK7onFuM9lVPlqXMVTFydbq9jLAkNXUgq+jHpfKLfumeNFV3l
mJp8YjPyuvuJAEaGdhVrYI0TVbzs7wr1voS/DDKIX3f/Me4DcD4KXOAw36zOY1CpvVC0qxBSPw9u
m57VIHdQOSppR3C+vtG1K3GFWhdrkhxtxX8gLFvJ7Ct/KMOsAHlaluNesq+B9xlIVUy2ZryM60tE
fUCfAaNjAjobOvXUlc6tq4AOvK2aQGdsfukg33uTmJ+hFeEaCT9lzI6alCbj4VVRKHn2uWpffgW5
yTEg9F/vkpn27hvB0PmTcKAAopXoMA0F/iLApVO2zsL20+up00fzwdhMtwfR7PdC0W8VFGS1Sg6c
QsVYyf3BMA+X3XqovMyAXH7IbeXjLsBCbKlVUh2gVvFKLUN+5bsbQ54SHdAtW9POdb0fI2tzs5xJ
YZeK3HlW3fzjMD8vQVbFf7sMXeGL8Rv+hXN5nYBSstoGyiFJvE7jhaHYCPinGATFJqgKIbm9uKrx
psOUFmd3y7kdWFXXTb9JoqUEBhVxFlP4sSWN0DIaaUDn0HE9Nfe4kpfg1i0JdNF83myw8uxsjJN/
xZcC2WbPQs6BDE2b8uy7VQjOZgjL0FsJrm0RUEVJ3WsrSpANxkOSNVfgd4orqXaU9Vj0iROY+uhM
uqe854eoiB808r68QjTcg5BN5DnevIRIs549wqyk0VGS5nHltlLhPGrNBcV2IXPq3Atn6aWe4W8D
wGXGu1av0dIm1M/zra5YnGJHbEN3m5ReTxfZEbyxHSdh+UGaReBHIA0ZiHN22MaBdcDYfUw6Ibn4
SvyPPb8ZIzSavwAqC1zi2Dq7cK3JkhYD3nfVFsP/jFID4IUyxp2XKeIcyJxCtxyO7BN11eJ7UyNC
23uyfYJc7UktZbwRS0AEirkNmIcibBIqgcPQrM4qMJ4EL6sRvweZsCQMYMFXItbcUf5yTnKAidZh
1KDVeRuGEPTIlOzNmlJNxSaOF9Cz5+0TVF2b8mkRI+v4fNrcgIIB6GMtQUgBCjJFW7uuR0TfV9BB
neoNe52QHG7Z4Nnnw0Yas75NmsLAXVJ8zfm1JACOE3tt5p6Wzcc2gaeRZd2Qr/SwldNta9axTiIq
fB/vEuVpe3BIlq3SQc1rXjuPA3o0BWWAXVOsn8B64Zgfk0wE12+9Jh/dMhbqRlvE5kncDKhWj+eE
QFRybV2Au3knO3Fow5yZHsjP+tTeuHkNFPNPT52riDIwRFnPjJiAbD6pMJZAc/Ba2k32FIQ+pQU1
4cE6MGmCZPmatS6TRBuMrAUd9DfMrJoeTJyLCMyOxuqRb6sQmJnptrb49A4y9ZWTaJ1qGErOQVyV
X12j2D7h1DSIhjE48latIkFUFhVc7+k2/cmwUvrFalzusVCDS9L+IfXT/FwCK0dhfAOIDX4lvuh0
iFI8FLugJWIZ4aK1lgrjqhIaxuTX43NON8+zLHQOr0mtEtn74BafLoUPekxGz9bCq5Id8RqJHcx3
bdFAzfEmBQjzVCgz2l2trhZktSgqV0qkbL1iPl+ZRg5CVZrDXyvzdC5FMrMnbbHDpOhVf95KL0xM
pIjKjJCNQDCysWlUsjlY6RGc6jwT9125ZNCpZUFQCYxk3yiDnNM1ucywYfeO8iVIq3f3o4A3Zglf
4+UYvQZuxQZ53YLYKP0aMdkv79SPhVn/Uk17gmwAhhe778V50dgvgUVkjlQQzXkh+cN3kelLflbc
yqfzlWRV0Ku+IUnkNhOLP8pcNaW04Dx5zPUxXHFYiF2H4jDPkTj9gm+QyGcAp8BUis1I3bGSMdx9
JKp3YqA/2Xw0Ar0Mc1PkHQ/OAWRm8wL9CnrT5P6NlnYP3rAWerutFqRz7jh2bMcalcBb/+fTcZ0P
iBZZPd9cmJanKmeFXp1tmD7ATwcEqOJLnumqTYjmAEbpD1CLM/eYBRGyg6eKzuzH7+z5yfzJ7Sn9
uhHiJtgp+0L70vY5QfZl6WstcBF/zyKDGXRXrYZwI72lHlRIvKIUEtvQPIvXSVS6v/P98iI99q3D
XHbMZfy29K4qZsTjYu/pQWykd4sQ4eLzMXv4rfGehk0BNa6d5NMTuqFZon9efNaaY9/sLQOfpQVM
g4bXy/9gMAFA99IPVWi6KeHC/rvDfLxXPqMGGAIPIWyxAzzgS4kROqcTYmaATEbaqdDh6EPi24Vy
LgCVO+NdOC2fuuEv7TCt5/1BNg4/TH+FbX5jBT0E6bp2hbLY4rYboSRDsJ5pduUiewLAItEwnunF
cbx2zl+b6QJ8gOdUkyhrRQVcRAtNNnfK0O91i/O8RxzBcyUT42P0iBFqeGaju1FfqpZ2GwmdE5FK
MD4NW3k/ypyfZHosQnu1tP0YZq9x8VRb18+3NQ3ZQDUGifoT7vOGKXQ4chfQw9wuuGNRY7JkFJA4
Z5vLIsrcf01dGKvNJJN0WTWo80qwck6WtZe/Vqod7sUW9kv5i0dru8pVbAiX6Tro9XxXb4XN7cnQ
Gr8682WIlZ5QMqUOTnQPockrsniCVgUH+PrcaUOvK+6XVzqXE3eXEiTzgTIPEBwJXJM8H/eonfcL
eSkunIYtT1n3ySA7NROX3CRGiIEsTgBQpd9tRaadC+Xc2OgifsUQ+CrqRPXMvbGmNqZel7rKiWRK
ZLk4WxuiJvDyXvK39HInfM+mfTAmBNS+wuyT31MCpPbygcvqLM44Zxr3d3R9MC2AeQTDZs1D8kDB
w/d7vvI9JdGAUYss8U6gUlbv07owPYakXw3P6eRVxK9B1n+enjrbD9E1/0BgG7B7ES2FJNfXz66K
fn2CVpBWKg7iNLwntFD6BXHDskaYm7/vJRzaQj5V6v6geR9VaPLU0AdnoqzBqlzlwSbzReYeEETu
LkujcjNezAvOw0iy+Yu5rN2ZfcL31/sxC9m3vdirH/gB5Ct3tSENr+NNbXGgyrpnKcxs1Rpiq1cQ
zAZIy43TUkn8oW6ocwkYlrP0GLUwtBaO7HDyfspWrkdmxIjEx3QgrIwSE6K/Iu1ezXuXx6FwWO0+
Uua1/n3Th2d4rnXTIoS/Et35C3hFD9R9087DDkVFlAAzXSnkZ2auj2A2MPLRyae5GFyKUw4P31eM
bhMThOezQulDKtqyMr4rUZHNPzANwfpwMlCA3T1fI1JchQAYlwt6h/4rcTcIswyhYEiqAMQ4/XRM
OVyzO69/sN3gNGImOIq+uPQ3IpRzgQHy6eqFCesVL2FKehIVGZYcckGvra7xPLoao5ElFuhrM+DM
qx6lSNPgV1KcNTD16l6R6dsy4/Q0uKyraM3iEiFFVVr9iqNDlNknQxnlU7NVkcD+11Aj6ONVFk4a
Sd84Rus1WZbxW8fxQjoWPPqBlpkVlwqGVlkPX6XpEVg10eZpMBpNP2NZ8wuddgNXDDvd8dlz/1dQ
U/Bd//3Zdn2AgMEZIfz/P9xkRXNFaZ88uTCba9oIPx4m6ACX0MqcihaXfsICZEdWugSaS8NvP3fi
m7vFUD076J8ko3GWVss5Fs/o3TvZ1p4xWAKa7/cETPuqHszZHxbUmQ2mq4BX5A3hWF2O1WozQPH/
2HvnGIktk9IdUM4ENbccpHsHaDSerzgolwbroTv/EXUYXKEAlPTUhJ8zDYjja7fLbkQPmbc/hDf5
XAl9hT+9WLazgQIceP7tYsAIsys/KLbuEPWgByb9Z/j+AYj6UOVVlpl6Cl4XuhGOYVD+QyeoKS2x
HSSrtBO/sryFYJG4LVyYslH++GrPgXDnLghtxPUZyXc/+NfVelbmTyDGhWkwhqGO5Est7cHScVgT
OOmfKMDloFl/DlBHyzpniyiZyQKqjo/nVYq8WGK8j+1pY5NJYiHPaYsxu/nGTNocu467trFWkl/l
yi/biRnQzaWls44RxLgVXfPnfRzPiPV3H/8OI+joP+JAmdqUALyYNctu4AdZrdM+SzYUI9Gx42+a
ahRlxrnrWi63VPfIFKDYQnS71S84SUD+vtiWtZ/29JZvmFBdkpVBqwaXPQUexg3JAAHxsAmw8R1j
jix5hl29NR9XnfGsSiFx0fUvtHnCwGqEXlyQbVL6+eIuedx+QTZgp+IZmcJk/Q3nk3SlOkC+E8kJ
kHyRaIlDKzpswqhIsAFhL+KseNSuD9FrVPK6b4s8++zb2goICG36fIww8XakSZtcqD9CfaGsOrky
fXzg2gt4SSKyUjyfHSPiq0HELtmRDHpSzzq0eNluJ1TpCbc8s9IVK9NEODAVxIKHe68pU9keSUxp
RRXLW9sk1rv+SSpo09yWxq8DsF3IqwJ+NoQJIgcnJW1UKiCxmQOcC/PufkDBD3FZZBgE9X1pdZLS
/dOm+hsu7GjQ5l9BcQHCRZFiYIiSqhDwrzxzFtTNaWji4pJLe2ieoqYc/VSdEED6g2vNnH7FG+oQ
kYeU7MJXgvqB1t8QLTffRDYdW8IzeisHp0enZ6D7kI7brcZJRj3/vW7wJtSipJFhvOtuCx2tvWs+
X5vT9zw38f1oip5x8UgzSvTs4PyCtuWE0XSsGtgrQMy30kkGZsIvXjc0I5U9WWoXRh+yjyJ9hrMJ
EqYa6DUzt8FPcLngWYoY977YSeZKb38FiCDCfpVLiZYnMz0EK0rxPj6AnnNHTOgTvLfGrrzGXw29
9sJ5+Au+0F+dd1ih7OEE3OIAPbDfMJApvtrN3PiXXaxTwcAHbZl9De0G6Vt4Du9ss3fSInu67fVi
Y3UxccXvjxoglvNVkjNarx8TrkDTehF7pelS0UVPgd7zyflmcxuEP85ch6em1wSKN+PNe6pFD6lh
VtqR8oxTmaR58NPvjacqdwLT36AlfrugveQiCdxQGKv/OaH60zZpHKjt5tO+KfKaERUpQ1Jb8mbM
X3r492Kk9Jo0posbPhrG8S/h5JpcXKX9WQQV2AjJFYSS65BXxdnSoYAYtYIZ3mrOCoa8qqQURj48
Hz5ZIJXGeCRZ1HOT8Df+LH4jl9dYLK8h1zHnZzEC5VafNfILHo49GeBjb1+yIz96JgVKOb9+NqRX
itMR/aE7xjcNDK2topO7tSBmSkeFehrRTiQak2lkAFsvkmvoNKX2++75waqC2xYwAgzSrk7+NPA9
5hpioJmiZWenzkKAJlXl+rLRPZLR73H9mrXmwt1ebYUTudkbaYjkB+lwx44wzUu7y3sNzEvdRVWR
vIODwO16gAc9lUh7duoEB8HgbdFiRyzvfNMWJMo5XXRQ8raZpI+UCmz3JLckePE4UO4tRrjVLoA5
/7Zcq5ZNxopJiMd0n1uZpWElLu47JdLIOb0oy9WWiPtriXs4TT1jIzWGBrBnql0I75wDfUtT4rtl
M37ud8KBOyrrP3XzS+mEmGSIVfRz3z8MvpdMoU2I8omxHB/PrJdHhn1wWbt3mgjHgoFlfxZtjCNw
tjhLzG6gU86R92gAaowOR0or9t3l8jgipyxlcsA3JtGsRxAlnvumGELedoTsH0RzDOfESjIQj070
YNY+swTUKulTiyo66yHF/DPno+yXrS3fTc538YJd8pUb/5Zr4wI1d4D5eVok0rHJ+GXAvoQisX5U
dVNO97Y9M+od9JfNySGDrIhZBlV/vh+8JS+O7rzUOULQsyJ8I8YeLsPZVXJN73eAMx07W7UfFiCk
Q2CmxCUfAt4K5/x1aaSKfgkkBlDF3gptAlYyLA1cabOceFIZ32JTknop3WrGejakFnq/spL7pVIE
rwZ1JuVGxkG+W7dzN6M8weTP1PD1uwWZDwou2bJfHpk77tWOQRf0Y0ecjqPSTS1C5o7+PEIAdkKX
Gb/mos6ZVLrAaF8+ZasBGzrLbVxIQ2mUVOl0NRcbQvD76bYAcKvyuj7mQBb3ODeeHb+NfjExN7wV
Y9zbz6ktgXjeC9hQlCGiG6Ylx+lo5HVLXyaDzGIGFxXjLQsHe1tyeAMmWH/AWm0OmdTmUgzV8GH/
QN75epPInFzVIz4YXAFqmDdOEOUVAvCCuWT15zB9IbVXxEknqqa9h3BD1OKTZfk2WxRwbbHero+c
z7g4stVPjN5N0j564hd0T9jM3Wwi+g0vd3Wx4bB3xSkZf/2mf4YzEGokaM6lYnwk+DyMjTBUyOgy
zqhrJONbpulFNMS5n+T+vDacDQnJ0hNjEHEj1Y0o6S7n65QaNB7HY0b8zYhTOlgBYq+X6jA5vv1r
JSLYWq6dL4zlicIcLJkqpNcFQo7FTr6LCfrxkyOo6IyEgmr6qAE+v0ADee049DV+SsV1vSUV1Uzw
E940ZoE4HVns507epInZJXZX0ywROORoSSxX9j8lV5nxoZVg53BBUc95KmpB994tsj9EPcuR8TNT
R7hPUrkxmQR3ZZhtEX2a/OwMaTvDRU4Rp5YPLxpwd+VuWk5go6biGPPr3htH+doPuYWWR/DobXaP
eayNjrE9aWJXeqnOIGKDRLtEd5Y5bT8CTGX5H2Ch35vZ/JzPmuwZHM5L8TTvmZS2QGtwM7p+u5hz
THUuDe0+THTuwleDTAtHnLDkdhv3GRMRYbv4RRAy4WKI91pSYxkTXEFXsOln7rLp3veFhpw3gmiL
TPrAg7HUSmGQvZ6C2lf8d657421lnOWgcHFjx45mP6Cnz8RFNnj+c9pfPh9C3RUb4Lo/PaQ9Dv2T
LNo/XLacfHKe6FFidnbMpnuVjx2tbcGTY5A+dUIrtYoU1PY4MZ48HXL8bFtQFFguAbm6Ux1mwmCC
Bd0tjfPfTR7Z/vmrrbvGbEucr/k81xCO/CKklbKsc5n9PW8u1VEr38lrH1Eqo6am5WwtxuH+4YSc
04AQCfPryjmWCIKBpcgkOVr7EX72F8mEXFhfku4SWgQ0J+O0SFni4jUdShY86nvM/5B7KYgYNGNf
F8uZ4V8zHcjE8r62hnjJfP11bDMcOe7FTWGwBnguSTXnjh6fJk3j0EUs2g9zS7pnf2utRm6No7ut
g3OM/9t7+j23jD7IHUzAxp/LDq7Pj+5QjLipWzRBQ+IGjzWb4GDgTzHH03n4MU7E7hdNxh55OwQv
vkwm0Vd8IQ7+xJjw/3HWrwqbGP8MVtuH1WaSmUGXnWQX6rA9DajOKmLQfPXtpezmNUtcpRNd2U28
wVEDvG7/kPxqKsSTF9C3oydCs1QA0LQ3X0JEjL5Tl3YifUXSCtsJRXEkTZnCIqVrkrdhVdxreR+P
2YDbdUGVDnEZGDrYUaTRp7DZg5krp3TrIO/cT3CV8iyi1dYer1yT4wiqPGlGQ1WpatZr47wzt9rX
+79/UgcF2Twic2uuCSvSBerClnQSz8ayGnLt7JT27C89BYNbiWKH0HfaOGJzaIUNFTDxE5N5XdwS
0HlQnuRatMNhhv0zp0dF5xmsp1QbWPkz3fwxcQzDWC6XPAgWeLVqOD/fRvrcqOqjkCqQJmdXmuSo
Tx69Lwd0mzQDDFRXIHk9z2etvSqPO/cFn8YZ81EIsT8MmoA3rpFoZ2Q5pFZueKrUBxPyp67u/R1S
HKW1Ti9e2iyDsnpVcs2wh/WJqP3lzCvWQi10nUmNDbujyLwnYWeOzP9aPixenS3/0r44KZdjEOYz
xbwoPjhM+oBQMGbnoY2WIVPzORfB6OddoUcRyrIqb555oBW+B5plvnZOXzH0jeIfC1dCQFuao2OC
9lYaplgc6THtBvpIQpcWCkmMfp2rv6WeTcswnce6gjn8GXVZuWf+pjRolQCsZM4AUGq5REGv3Orw
YQtmHejQClcmKfHHiPztBQaiYlXYAha6nEjPR/7eCdiKfzhC42KnQYut5lvU1hvkSIoDGG4gm/Kx
iaml95REvfG/e1s2FqZ138DqxYTmMHEAWnbajk0b2qTdETrCWaXwUXHQpzNPFSbMzXUuyFzTVioK
VeelUSLki0vprKKEuwvYmyzfpXO4wgOcsdgPfy0jlhwRQz586mPu4fjUF7rJDd534+CdkrjVqzHD
AmUWU8rMFIDbXJZrNZTnR7VwWgwO6Lq/uV0T8Pq3whGgb2CKhw/1BvQ1D8+n6G5SaGuZSUtjrlWm
fGYunLHB/SM+2NlQv+oRXsCMh2YMDaVr1IXLY9KluV0Hcc0vF3vJZOPXc2cq+xF+6s+ZRRqvZLXw
Tc9dKFOHCe4KiOj+wNIkdGsn6e1J0X1gVFZaGcNFuEYP0SadtY2RxV4IOQSAbgkB5Hzvn7Y7RFYh
8uYuUljP9OT94OSDhY3896X/1fla2v3TUIDeheCdn1pWNK+diJ+bumrT2wuK08FbMQ51k6fL8mCG
WcM+Mnf9rDrx/DnE1QZTt477M1YOmDO7Tpww0YlNa9OiVAaLvqXHbopBDR7HKprHKG6g3oUoDtFy
ty0f/e1u07w6jg52RrDrqWGre1Yxl+l9bbj0McNSM61NdEUi2tkvLRA8svdl43LDWxDz5i6j7MCt
mSIGNaQnAaQ8VvAJcza+MU112tORBNOPfGxlwmxJ11EEbZwtdg+1fWStFjt9fv3RqclLh5sM/Qx8
NRzNObw8BNvgtKvpGwu2ClWt2/HvfW79MuJzXSnReNptPz7g94z9/pzWREDWiFIX/+xjvX1TP+tq
b405SJo8nVq71QrDVi5MhIMlT4kS1ibLGAPybZmTe/PF/+Pq4ZY5RRzN4BdoYcTLCvaHbtNVHhB3
p6La7Pq7F4HRBu7/Kp8Or4HFFUMq/Kx0ELTQkI2k0WqsEnXIo8pYxZlXIJEgi98sDDjrAZFOE4B7
NkD5pE/hWrYrMSEvizHlJYaj25+vIqx4HGKZoI9Qr2dUuwXitRht9rEtx/VwctNG4s0IeWACF5UZ
sXN2VE9O+H0w1clF1L27LT0KlersLwjhYZq5kPzu99L+/IvwWFZFnre+V7akmOzbsf82+qIZMhbo
1Ktbt1pBR5U+pBYeh+ITWla5uH8bq2ulsznBcTNZKhhLP0zQPRUc3UiPhZhdEu3ZfMoZ1OB+xdtg
vMzM001n4htjp8RKLyjVEvlG7llhpFRCYYaKBHHGKe0eJ/YqGMsldINO+T3A0Kl8/4/PigdrTBmh
Q5MuyBzZxx2jPBinlc++p0H/oK+8YwwDi4sJUhS1fueWJGoj3IXOAWfG9pAzCVV6MX81iFRh81sr
FDLM5vnW8pGxcLL/ivaBc0byHX1OlqVzT5q4+1IiLLu7DgiVts2qr2DvhV2rkX1VNSnQ+FB/zoXZ
+QHlHD/OzV2yUQ7e8KQUMGmdrpUCxLYT9bpR/qxlxEYioHk/mGgycgxCi2ZVNfnYCteoLKc4iT+u
HlFCfa+aLBw0Hle2POvBGbTH0O86HjGMEp+jU1zb4YmzTKgOzNRNRdXxd+uYqXI759BxwrshszKv
WBFQ81VESWqvp8V5Ajyf43TcNQkNfII3MoTrWboB2yhWa8HPQYQtFofJ2MP1iLIgA9SyI3ThI2Ks
feoNmG4K8cg7sZ2WNam8lCJrH7gUz6IFuG8PTxT74Qu6DKFzft+PutCPG2wG/GFte4F8ZgwcCDft
yHdHa0xIiOMWNJYDeOJ15KNG1kqWmBjomVCG2lixkTh0VOz0zPqGBFT/J2eu9h6u9fce88JJ8Tdd
kPC8g4uEiPbIucxfGGxn3F04idqdrPaPI/xw/j4fhMdXhPiKzJ1agQg95RP5N5Jniixs9OQfmai7
5Xo1E/uIQLs5pHAZAcI4N6Q8GCy8m0ydqHRkUB+QP4vQ0EYw3HOl51uV9ZVvgIPJqPnMAnmMwnOd
iEUVlqc9H0/etfoQW//ayR0e9g7peXo3pIyG2plsk/GiamkOvMGpfjugM6fEwuQA7+kKnC5Ilcov
2S5M/JkjScolU5l+HvfYSfm7ojbaFPXjOR1mR6ALH8t54lVz88xlNkDa2PGv5Pc8Q88ZIa+QDP3k
5D4tn1KbqI1RnGUrTzx1l8MIUrZMmxvRHULzd1xnq9iUEz+kJa7c+P9o2p/vyNLzHOZrf//g87JI
qBuosE5yLh04vn6bpX4A8dqQxz9EmNVFD++8mABD5DhkLHI/ninz6oRZ8a65gfuuH6Wan4rJjk44
tUujHDApNglHh/bp0WfVR1uqoTze/J6jEs6Buk0JylxxD6pox8tgnQjjw215njYhJCx4t6ND9E2B
+WSOgV91brrWhBfXYwn3hACUPPj1xbayfUkR6FlxN8/bU7WnBdPtAO3lGNKtxJKSQL1Z6p1xTJb4
lz9RHoJKQS7CZArWEVwVLGDG7Mru64ZYq29rvN2issyHvvQzjc53g1Qj2eCwCsXCr1zlBlSfVv3q
HGibv7EIFnf3vbTVokwcswkKhNrP15UJfFegf/mriVG8AQsIJ4XN4EoVOHoqqpbAoJIbWk+wQuWR
GqJ4rHY8wGIhvuD4FvUF8BI42V3caG1tDz2Mxp++a+FKySvX+eMfRcuW3qIxsMeS2v/1PNAHVNKU
dt4LX65bx68g8o/LOOVIM2nVJ7HUK/2CNwY6tn0QNlPQOlSQiquONwjfsNmmyXfHHsp45KJ03IiO
9XGB8+nLcxMcXb4+g9q8ogOnMaxbIVAUmiT0ssU7Kr8Z/3lThK9Gisg07UKW00nXmfU6Oo7+6X0u
DU6j5D3wgmEd86FnZ4nywK2+Xo5d69y+k/ZrtowfN9lJ2PADA+W+vVrsv8lyP2WPXMEpdV3erydw
eumJu17PrGTRTK7EZvobxIF4O1pChGW4iJheDC3um1Sh+/VZ3zO7IOAnQtkUtjfcEAe7hPEEDuTF
qREM1xcjg0Mhni0rQXHhnzrRWPSFjD+5/nlqzHQr0Zw1IWZvWTNCSwZjJfzVojvjh+pFeqtK18af
oT0MiKvP7+2XyEqI+mS4BiARd8fMPRbfVBOEulPPOxh6wRWzVbJlnHHgTbLTgQCCIp6MQC6BNKp5
RDuTcULPD2csBav4NhaHtOrxNnz0rAPQt20tcOmRA9FPnFm1zctcv5llD4cpxyG2JuqfEMD4IoVZ
4E90jzBVsCoHWkzNPLlbo4T43NSxf43yLr58dNtb2Tdc01cB+loTUEzPnp4o5hNg3geJHuluhrM9
Retjs6/9p2mxHSPQmC8bMLj6NnIiU6rFaBuGyz1U48Ik2hh6HcvsKp8aj4dDTRZTT55/sPJNwT6W
RPr0NTEzgHSfOHF0U5zqgznDz+Jg86EF3+fyOQF18IDULW1DfM/h30/yUQNI4s4TtTWvNPL9qGui
HjLgnDnEBcAzSuO4m8kAYXSH0l0IU+/IXn9vGhG7nvkOwvms11CgGCAbMJSue7nQxjBQKAWN9I3z
rWTkDoXO8Tqst+wXnm1jrtjE1k1hiQ2XPn3zWEXgdeISnQ5RlnaQ3X9jSCiBA+88DIBonlL9rw2k
AdZNL7/gZu0toE3GNy5VPL47eED6JtXM7scbnK85r3fca9h+9TB1u/CO7wOcTZuaUcAAVldEsBvc
Vtc0dCMgC6xBW4muvMdViUSAVtwFX1PrgPbgX7ldc+T9cNz8VJdhOJV4Fu0gSjDCyf8wBhKSuJJa
1JNCGgz3S8rluxV4FH9wV8sunFH26ZOJNvBvsB/Hphm8LwXhTgnzCVZJJJAa3B7WFlSkzUVXrP18
E9mE/Qd3wFgurZtFxna9doY9ssIrUda7Btq6OIDb45OsYq1ZM2xyauTJoDcn8tmssstUBM8otIOP
l95hkIhux+K9ZXabnkIjHxeHwuu727R8PNce+nY/+lhiDHVuYKO7PGLbkDcSspWtM5Mr+jE2r0RN
mQlwOyzKjzbjxVxaI5ZtT3A3IKaVtiiGJnJTv0utpt5AaS+mfAVZmFs4CHmLBYGDZx/W1NXB058C
q8kKNwEpGPahPGfzfHe1AjdmLRVFNt07T/BhlfYT/FDbyasP8UhEO93Y6xARiIYt+r7A+o190OfS
v7ISmdtn4eh0SEc6vJqH9Tg7zcBU7qHtbD68h4Md1Vd/7WI2ynHQ0ATx+zjVMKzRvDwxX9+oMDzB
Zx74csI2aODFBVVrqPnCady9zZLEUF4otVdamzO+HR3lGb1NcSxSw1G0uNqeJhFEa2UdtAk6jqSW
4kbcBFmQaoZFgyKLMqNOCJnNc8KBdlqQb3RRyI+7duPOYUxriSPtMFl7zAtte1xXs1TuSiNIyqU1
2e6uz1mh100jGC389MDitObR8idQ37r48BQQQL75g4YW7CA2uokvUqhDLLQ6f6HFJoU5FXtQiDL8
LG5xZCC0nFcyBW6CemCCWqB2R+SfO51/fBeWAgHQAZqivJbvses/rIV59jL0jfNA3lUwmmDz4yBJ
RmWuaAvw1P3r6Y2zh5XTMLfiRWYijghwB1iLIL+DEud2b1SsFbPikJajTCmLIiDhIupH0govmJ/C
7Yoyg2lCxFWwDLwtqgbUt8mWcUOlMTr+JOii0ImmoCDOekZ1k784eQAtzmSwbCHZhmc9xyQ7tbus
M7RlqLooGSHgbNxNjiRdy1wgVtd80+LcnQ0bbNIrFfJbtT0F42VEF8talG2kQjfJ6G6IABuMl7gn
N9qnA304vBKK9+wrm/dO6/uiSV0J4WIpe5HfnPjp7u054TZwBZE/1drRjoUHTlaV3Z/IobNRPNIS
XS/wYQDA93NRMxTl+8hHt3Pd3YUKyA+0BdIGbu5V9Mdwa9LY/M++oK88XMFa8MgEePsqqloqmvhv
BaqqaWFyp54pQqPODJASvezodU7on6oWQCC34OZLHuS9KLem/3st7rxJvU2VNd83pHaOeZb0oFhG
2oTS1fhrQvSY6FGWoTs/NtKu3/8kA3rnKeQhY9FGhqs++YmP6nkUaTKtVcfiN8M4cZmC837KiIAH
rtEh7xP9Z3JhgELbz6ZKC9DuER42io6trTuFd6ZIC+BIQLCs8bSbvLfUcy8N7G4dFeuAn3oBrmHs
aZwoPeHaSCpyHaIMUHVusU2Zcaf4cf7xwEvDHeGDrUU6+ophInVDr1bzvTJLqt4yTxFxmVLKa2+t
GYQWPhoOzEJSiOrD8d8z20n6pkfgWNppxJV05d3DzUICf5dTOqTa3mMva8rOJ2B18/LfJ104ec0s
7HUVmYJIcb4C269uIw/FASreTYvtBAYtqAsXmABlE6wx6gjHvyEz+R3fnEuID3n8BZVBp12e4cQK
tdlpo+tCJgfTb0UtVtu6qHfsHBnZF/NBSLSkbsM2wCjqufpV6JEutYTpqrsHzHyZWOGRDYLxxTye
uUWuV2PgPRI+k6n0QBXHuSOIR65RKYJnh+pHhod1d+5PlosVGZTV1wzVdUYd7qX8/+hYKlydK1xF
tX9YjXUwrX5wfWgqnxA2Mtep+uhR11FyThz2SrgnKaSdZoO3ODHfFqyBpBqidtvVBcte1OwLsBLY
F/fdu9f1BuGgBk6aC3SIE5FGwybh8yFwrUzjQp9bq/gSzoNLlpZxIZQG35daB0SjQp7E+RIpeaTo
JtRkAPmz9PqM8tEdg/AgSptSRjI4hOckOyP8nTTqQEMXtnNNnX3ZHa324OZ2bQ2YWA2CshOIIPfE
B44g0kHiDOnUC5gbdwIKuX3BPsSDsLLB+7ew+w1/R7pxbYB/yAEGGfhWbKz0FjzkZfbN2Zd/Goxs
LnhsJjEABPM46BeiiTHvs5Cj8lmtSjX63d6pnogBTdQuJv9Uxw+h8sAvCeioul4Hhv39g4eGyx4K
ozqGkluQWQkP+Re6iyVSorfa2EyXKt0LfS8Pi2Diyb/KCDWuudV4nK4QpmcUJnvubQgnjMw9v2qV
oaaMMLfUoLpSxGr+d+VITtk5rii2jeF6j2jQMHMeb0n64ekmOXLLoMcZD34RJ4YWgPEo3y+qSgYk
WYSJfC2f+NqKMePT3PVntSPZoAzxzm2/tX/ctLD8LfTK/o3oWMRQMCwyrFQSaoMTkME/zcfsRXTF
Wf/JgKC1BDW7EDwqw56MDugbSNAtLRKEPdwA/GMpZJbm3dyfRqGJen7U5JBVVUMyN75urz3LktU3
MDBXmxduFgcmXpeba3D3lZquMNk99HkzNLYNxoeAhbFhpZN9Wb7Rxj3PdmaD4GP3sse4lfU8VJlL
wkilgBgd/oAxC/Ma2CEQX/ANOGN0vYh+tIjczjfFzEP1KhjPBczjiNY4oVe5H2Gp4XMwAKq+O8WG
McccycyLkMC4Ru2gBZ1utuSHPlj54UckbHjw3+Txs6YmTnNMSaj6TOqtqK3kar2ZKqaSpXZvBdDh
uOw7vz+7I5TwiGyfgAu+Gq26C+6O7joBmuCK8wybMNDYoA9jjk25fSpbG7gngd2NaUAs2XWE7iKm
P8n5pcW5wkehGq6VLmWT7ffX7XNr+aznFL7P+LxV3VcV2ZMSZNc9cFytbGO/UWlbtez1A7V1BR/C
e3/sNRaUu2j/EakkrF5mj8t/73LWkJWrkKQiYB8orReqi5xT07mdNLKJLUCMrT5hkkkPFT+6bRR4
VoE7bKAWX/jwB+FlV1X2UIzNsgKy49rP3fpq2C7lxnpOy+ZGehbuDBhQzoqexMei2Ia+6vR2OxkL
oUabIxGeXyR9mLE3aeRdSszYQXMlL07/N724OH7hZ+H985yTu13rvkfrLYIMxTcQBYNsz2MIjfnq
4+zay7aHBUzOMrpPuzPXsK2D5kp7uJiqOe/sjp+7sFTqkfTuoWA/Opn/671ogGTHlbDlf1v/GcqL
jxHZ4Mvfb6rhqdWUQHZNkmUrvFDgLFXMC2+Pxi00LDZbjKmD7i9+CmUJB9D3Qy0KN/ou+5El3mYn
Sc0RFkyUW1dc5ow2qRrrvmnV5hs8LJ0hyvsJosVWMl0etocGrwQ8FOq/7FrRudKftaIdhI//l8P3
TzQf3vJ3tFlTMGh0YsBEsc4SASks+OnMXRm/NAjXa4aWdB0Sg/Ic+xTsuL0Alh4417Zn2vkzP0sQ
ueyUVreacSz4lv58P7kBkYnrx0Noz97F/25tkSNYo/0YHQeoGZy+LS1qHozZA64Aggt9Yl+NDdFY
XsGczHh4akiP8aUgmWRSWxx0+2n7N+bEArRf8tdG7FC/Qw6+Ohm7ljWY9PyKN0tuE7uxlobdjqcP
4iM3cD8JiPn3OAd+3J3q3Kd2PWZMHjn8i7naE97T3qfqfxhSdbtkshg0FMlUZ3hDg5DirzSCk7UR
459E/U1mKy7F77w7FJ8zc1YZUTYYTdjnrAGbt1xKcYy+DeFTRJKD1E4ZJKBPMSvKbTqa/M2WE3FK
NkdQ4YuSt/K4TG/BTzG+K0l/jX36BxWFEPH8qBff6qvx/pdasWJ8wjxG78hHocHGX5oxv2JcoWGV
xPlT/dtgSBZLGW12OY1/cg88cDZI6YNGrq+JBOiHtL2oCVPWm8R+5zjnXToMuY7E9fKe82d7NHDA
pphx6v8RF0kf8D4vSTPSTrRTSowCHGPyuZHmAa7V8+5Fb0k0OOY4GO2Z7kmfz+W3X3r9jfy7yjXA
4flSj61XWJ0vT0Ebpi+0fjnsLMX21khCOaodPt9FFPHfHfoZz2fWlUy1Csfxb0SiBGNUTSg/iI+Y
wCmfrzSres/bLSONsgzWsGG9LRbHrJ9vvvL4PIL2C5KpqQPKJujYbS2IuyFMJJkNjuTd8YtJnrjW
H/YGMPLqxwo+F7Va/rIiwkR8Ao1uXvS2cGr9Rfk0vaZhxf5SDUqkGICV2ST5PXBftuERNDQU10MA
wld2DYZxMgOOHLWj05c1wboiNYrG16wplzj5iN16FWRZdhHhj4/vC30rxDDew3nBUcEcaNNPQIzs
FP/ANgk42OBIwI++Se3bU3HEbBOUw+yVFH4bcqKbpvgy9VBQkUPNGSEVseCHS9NjVnAyY2nVT8GA
7iybMxOu3eul8sPNPZbTEstx6lXtOsD5Nm8v1bW/VqIIg6CTctNyVAwNrPuHq1z8jATvG+qKWNZS
dgsIiEtTn0gGf0BLyOhhKz2LhyoLCmezTa2tYv+PaIbOeui0dN/ixWJJz83AQU/woTtluFmJdxQO
2vldaGUGcTBhbfAlORS09e0CzQcdYM2QeaPbqazPHkr0TLiyvyqd9D+YNSet2RJ4wcTfz0FlEmh9
yCXEqRCht3iTbApNE8P5pBEEWZ8l6JnkGooq/Sif3aGqYjZQuZHpvFiGZSSp2Xwmw7X58aUCHXcZ
RhZbyxOdQwdkn/Z2DA25SoS41V+QxOYI2Lsn7D4IaV2ElmJYP8yCc3hmx4Utk9/7xD2jYXF9ZKMx
NpNZ8Z79JOo7vzp/WByM3KGAi6IK53C1eFm6K/9VF0KP07vC1Ou+N0R4Q4montHGrhlM+sVs2Xll
v+S+NF6vjW5SQwytHBfESauqzf0cZS3d2I8S4E1OF+kb8uXW/sRAKWrk4Zspw/7z+B4halVfZXJh
32hxu84+9oMhfFKqigDrOBN5qXp4JD6zNEfHs+HfG+Ynb12D9ABhlTZZ2OXDHBvmFTchzjTLh8kt
qnK48fV/M89bCZiMB0eXNPzDLO6/HXHr2UmcW074cNfP1z47oq+niIge1Zwk5cGjUZAz/PAbIeJx
jysQ/yO1jYjWfHRm4ON6uzJkCMvVeeOo1ps2mS3OWe0nAyNGnJexb+qddjGKWhcfMcvpl8xZE/re
BMtMWZcEDLZf3WSGnKFyTw/MadRnVK/AVMBkaUIkD7LU25VDW5yqBChJ+/p2noekw5/uPvFrpYOK
hrnmKWeqc1FrfOELHEeEDMYYBwNG6ZgYGlBazzVuQR80WbcMwLkk39v3nittXs0DNw8Ab/jU9qAc
h7vWNHEQ5L+pixovnbvb5QTJ/2eAt8A4ISQZwy/Q68sUU3p59sq+6R/pPKThx8MFuh57BLzkLFoD
DVQgqQIHI5yzr8bo4jzqBHzslNxM0yn16db+eLHbKCAaHPJSEIVkkZssGUFKBL8Fbtx4eyLwYUCK
Xcc7iUwuQXDFnifj6XQ6O+9noIqyPFE5/M7DMiQKVXiTp9AMxFUeln+wxEB0l676fBXS8RhwTDzK
GYHPX8Y/wG3zeLbLj1cceuKVPCd08ts3hBwn+xqZlefatZKgil+S4Ij3FKxGw2jsPvyGvQOqxpMD
fiAPLTvLjvpIYuPubtzA8dehv06ByXcz4TM5bVXn7PvWk35tqUcQgHq8bKRvEl2Nh4g10hJBCqdt
8EmGFwNC52oo8pPPwV1REePw30UaPbFaDGaVsGDmDcY+KfAjEeIox1Ir8KMP9cpFimDYts1F8qeC
i8zbiF/CUNHaHJKMtjHx/vFBiBcfprUArSnEM/deEF0u3XVQa0zznEHBzAd8OeWKQWELVFx2nyZJ
iPOo0TnUriFXG+KX+QzRooKKsspJRFh1zCwaqozBjCBU7M5yERRpEvA370jc2yxvphC2w0/yY8Yn
sGYORtWu0DKkjJUhje/EXQ1wJixUov59UY0seaEySAzxjSvjzUuQM7Cn/DtOjhsvHsvCvDPq9S5E
xPA/2y8jfQH0cl3gFtwAwUttaZXfdhfQ9/djwBiJ7ouHk7MVZcz5+Y51WEqoVFC1wQbsY2UMd+0C
M1ckBugZ8B9P7pvJsYf0h6Dl6k9/uk6cXwgSkI6gnMwCP8wq7RWcnAbTwyTrp8Y8tpcbGE9sfN/K
engcfjHVp0sDNQnlJ5C+WgEL8ErG96pPb7K8HUFMrVvNczpyhkUEZaiFEfuyHhXnv9hVwtEuHPBN
CJdELVHzFD9K9sIlUOFY5tPqzwMUeoVAZTG3/4KjufpQtbxR5JZMJf02MBFgPoPkmrdnd1ZlET4V
oxlB1N7+Rev9cfamJNlG71onuNW2b75BVEg0WJOMfGa4DSRmzJCWk2UxHGN0lWkyWFzS0L/LJpnE
TJNfxaULgAh+EUbf+9k5xFHBxQphhQOvo8wQ08HF5hDUbtpjEB096FbuFzY3GDq0oEZ6cyfSyGjG
r6HTt5FnnAt7L3bc2D59uRlqdql7+f8ie5QiN6BU2DtnxXXBcP4kMrP5vNVn7GLZ6ubpuAtf7MKQ
sLsWCbKjkb2+WbnzKnx1UL/BqqwIRkRu3jxWzNMJquqk8mtmloHvja+dnjAHbZ8gMXxRsIbyDinN
ezQXN9c6bhmm9cDDgR3k7YrLGE0BM8sUWOtd4BKjQWerELYLfkficcnggEyELn0sHXlBx+LPYO3U
K0u0yg3fcrCYFdPosaj9KeYXzhNJRk4l3Fs1+Hq9dtgk4tTlnRDVEfLJ5JmQInY+5Ap/ie17hztv
+OIoGP8O2XlJ2EBZARn9a91sOueyAoJARmRGgW6AmAu7L4jIL7NjuBWVr7XYXhgMY4ERvoPN1UNy
VMvI3D8CzaoVv4/1Yb9MkSA8S1WWKMGgHgQlMhxpegzlkeGArJr6b8Rri1x6N/X8BEXhLUyFl6qc
gq2+yPu/heNGddFCin949gkM0tntm4VqPpD63geaKUwf6sX/lA1s5hnpaRVMpB0axfKH3o+SP1af
04mHBSNHY9ud3BIl3eqs2fq5ocsBX8URtR8lOuEpP4/xkOYPk3ngmy7zUyNmpOpgWFWgqa5znfx6
ueGv2B9d37i7JPc3eSyeMR3YcQ28zVU516WtgFHKIg7A6km7h1sSWK1bWdSQwrVhoygfnYv8jSAo
zPvVLS95XPZwPUN8lThveu+0EunTnCipCd3645vOZOfdDFu8UTmWHKpJW6Kci88gbn/HlAsfjKvt
7vn2afHyV9oRoxSZXNVBjtQk+9n5LTQbUxEW4cPVoS0Kmsz/Zo2w+HFCidv+DAwuBvJuC2kVrD/W
H6elblKYfRrpkwc39Z8E2fyY+jZRAN5lc4/po0b+exr09TAJAl3xMQktXziybcsMZLCNadyQA3So
x2f9VNmjI9N1j4g5PdiQt6LViPJSYC4CE33fcjpmIR4ni7P/x2OjuXX3+oQafaZ9RhtcsWiDgM+z
cwACav/lBMGMlHf4OTihaYXujMQy5TrhnbfKyHqQAyonv0f1+IosapAZuARQ+dzU4LfQp5W6ZHk1
joWQCzEqyLGTym/tjYYmetfpoSzMLtpBDBJVDQIqneDnKKwx0ImthYqKUzBU4Mcxn+kqWREvJcz6
ONjYRPh0iGI4hKZ5KUiUkAthwGuZB+ISZ/a0htgt6w+BS5Wf8f1NFK/ve/1EiJZ+CvkXsZhzeuXj
dM5yckcGWg+i0WU1B2gKbXij8ViFY2iHByz+D8pn1z0oincnw9IjG0q2GcoQj16KtxGS6Bhg2TvB
CBaKByQYpii7jrauz52OOIryea2m0BGhrnjdIsE83utQr44vGHFL4Zmgfqa6zEc5uBgEKLlKCbFM
fS1qAtdSGPdCn+H8pUHskgHBFnytebQOeAHHgASr79nBI4bMYCBDsh0QUddS8f16jXM/+2OJ0ij3
sKkwR5fLolN4Gc58jCOcA/NTUFlAdhwH/b6WHjRB6ZalFriYASP0uvS1oKwQOW2Z0iG235igpVn1
GgtOA8xkoLtK0BWqCRwg+pesMrPL+4yePnF0gEnfcdtcvTXZVJNFwTFmA6Hliv/eidLHf4PaMALm
uA7j32fTUzoof1IO8DNguYfcDcdagTDyzvvXEtyCAE1YLeZL4MyjUq42lXtHsOGDOQKzRQA5En0+
21VDJ8rY1VVbsVZ+kVFpEeSv1gx5clPf7lt1RlisEF7/j+s4M+DwM1oww8Ba1/GfCBZ78+Bp8y8D
5mcObtSDHQoH/MaM4eypIlUdIQBqUtdtuzjJsioE8Qpwk+8e2MQqGlqY47sNSh5PRPuz0T9cIgdU
UGhVBALzzsO6TcbRa/TpVsVf55+TsB8wowklVSwSsoA1lxRJhHR6Y/hbnVM1h5veN50Vxdzn1iTp
Ye4PaZSQL1F2KIQA2JM2CAkLHHK/9Wxn8M7fodZ4jfW+e17Xi88PM28nmKXuau2j0XB30n+AbAEa
O72WS0WDX7U3K7vQlkcBMt6RYxwnwBqu+Rrr/9GBxfM+xhkGe+zfFtRr/ctQm+t/MGqFgCL219Lz
1wdvs1yseewS/cOFv2Oi1N1CvbG2sySGIo2X+Pnjdw4yhTxJNmRCyWwR4Z2e4cWrePziWCDePtYc
oh0mtQ/FXYGufoJBdmzRoUDnzNDfB83Ppf9kzDNRfn4y/Mx9DNoF/PeYA9ZztJWhoy7JN6A2dxNm
GdImu73caU2/fYhuWjVPv2Cab1Yyb+P5I2EssmZ8OchfS3lAPzzP2tDMwUedqf+MLDFRjJ9g62UA
Dplt/8+l71pt1Y3uecwVwi+QGh56fduGFRqhbba3CmcbcuwJplZVF5e3TgF794xz22LL5WAa0Qsp
o6XCD9/R+FVRQazpAW4rnqZlLLfdJPw/N4CrhMqlsmTpaR5JR83fASs0QCH1F0vynHgGvDBDkw5D
4zgvRAgpbGrBVnzgZG6WwsYmeBWNAv6v4cQ6MLJMCzNzJfZw7qcDThwndD04G5RiEPsuVVyoq0Tn
9yw4cReio0mOgEPhyad7qQDwotg6Siaa2VIFu7SKeCPPCiIydqSWDcnsco9qnYGzX14sD/tdzZyJ
iJJBUHVKOvoXsitpKqLVbRpOvSDYisQAhTD5P58i0kjpfn8hxDHKynXFCAG2kTn34hOP1viRi9eV
PcoOKpTNBPSeyaCGzvUx11I0A0M8FV2rPkUmP+uhSNQzrnhbcgYdj1VhOfDUeXQGguFJRpNzIj21
aRwpFTkBKfTBQ/FWOR91eOe0sSnqqZKb8UD2xUP4F2N2ws7fGGRkhJqXw1Aw1dwTvfa2M0rCDLDp
UsX10P1SKxenb8pfL2UsYhWJsN1TEvW3cFU7tyKCjPwj8sbz7QKLGSazpd/KLa8bbLanoTLnPCT8
HKbcO1blSk8RbQQhAnaCI9bGza6qP5KDGniysDwd+1vRKy6J1U912Yll/oY+GbpaR1w6S4UIb8ZS
LjIOZcOyNH//VqhzZGBPzc3s/gCLF3Xnx2CpIXFxRqpqf0HKHshZ4nr55KI6+a0yAhUwJEosHNiz
bTqOfeqMYbRCnnAzui1BhrYeUu8QdcIe8pZAxLvEaTaUgk7MEEn7AqDH9ZsKT3gr9V7hQs3+2aaI
jpxvcjLyPykMAVWSGCd8RVcaassPpMDugfyctoxxHPoxfJG3FGLajo8KKiZ3vSvIfd8m5yafDKpP
K9tLMnsXROKDbZp+N6rjOEpCiKA7DINdBMm9fb2xv3BwK91mukNyYBnCOVNQr3Z0LNR9Ek8490ZH
KkQQVSIxcUIsrdMwDLK5xNFqk6hTu9N2xbfWFUkwOmPiTGyv7lIyZy8F8+GyMJQNZ1VZF5RbxRbo
3uLltUZ3rCkOSMdFxVvnuWJRBc5QGeLU6TiMNXGQs3GEssxvePr4brEbH5dbfq1Va2ZbI7yABjQF
t2l2ks2jSM9k3BOKUrXTJbDIgIYP8TY4oei8iOciTC6RtFEQkHCPXN2xdDdaw6Q6mrHjQwn9Hjwo
CaDf10LUyAUOeg6O2+CZYAhwqPr/iZ4Bb8Hq5KAkCDnkHz/a47SMwzMKP+yNuW/5pIwtScIBPQi/
sTTrecu7nlIGcLom9sQG4es2c7OoBHraNcN8eFS/UABUA6gwYzAQfO/MP8WF3JrQsjaebqrSNrM5
Ojvdi0+3NeNrV8qygGwppczaRUb7lKOVVjgzyW1QVPHMju8Ic8U2tRXI5qNtTAsQBwvWrXkVbSoy
/5T+8lYVQtmC2OuW/05ovBsU5665mlWlgAwGTSgVFAUJkFPgrwQN4JPVybqlcYPgl4quYlJn6LhO
hd1o/XqRWEP55OjVgDC6Q3ALfMS3PWWDhufqjVe0SP8mPDf3qBHpZQSR9J2Ft4x7RpTJWZgHNu1z
LyMXaqcCXJXrI5jMk2S2JFAkmUXI8QfHerVbup1FE8td3bFEHot/t/X/0h1n7n13MT/B9DM3uVHE
GP2TOvEavjTkhU8ZIh3zVJShzRIUwYwrdRGiUmBdjOoBoUEZGxqIUaN3itDrSQVobj+DRHtZv1w5
IN+dY/JegmF9tOaAjo9fbyd5mLxoW/9lvNN+sLOrdCem7fWo6gjZA+Z1uuEVLSiK+okHkmmRp0n9
DZMGP3KL7Jef8N8TEtNQPsp6uelVhU1n0bS5WrNyOvzZ5MbFl+SjYBr002ZKx4SIDo0wYG/TeQp9
1Epz9tHCVyyj6YnehDAhFWjPRM12+TfiMkRvGXA6EQr7EyBG9cozKeGmqD9MmfzJB4HZEh/TWYon
3C/c8lCbN9vGL1UppUICTwuX9nxzv+vTbep0p7gNW94XXPrgLiwaoohNFbSJHAZqf4coxPnwrBrh
BOHk1AbH5kpJY7eeuqEA6514ilPHaB9wfLa+/EaOTJrbqN36zCv5bVx2PT60fSWk34KVRFcKKpuQ
uk27QsRyJN/uDi/AAFRB0n67jQX5G/SClIPRSS1WhjfkFwzO0N/qZPwrlq7MzJu11ZqfDau6SoHu
mxT9pA56sFRQ/tQyl8zGJZU300zXNQxBLjFpwr+BMXgTVQ7mHZLTKdAxlfE0IgsTziiVvvnaa7px
Z00P3mQVeokTkFkoM8QmCnBX0jxarAoRqfECBcTuhWHzwaZ82KHDiZ/apvFdKJAlLBoaQqd/DQqk
pcA/TUq9rzWcGQz72oUEyIIxokN3/uZpMmyBxv4yYqcdr+cVltbUB8vQ91p45pvCTZn3EtB8MhjH
ddiGMc45mC6umgY3Ku3qCaeWi4XlUqU+wyF3E60nRWL1549bL1WBw1HDwvB1Y5FpfcSd32/wVBgO
xdcLqIwRDw0RvUX2PWLeaxw5j1HSdW0KUKUyeMMAOF+tPuuhnkLsubJu2dQrDUcUjVoI5MfMA5jp
cDyXhd/iBCmq3NdXXZoMFwmDjNaurLSFYQesjoFYAGOioo/a51gQQSWbmkhbMU06fxbcBN+4QWaP
3Nd9l3O+37BnRcdnUJxXkmZtnrZ+ByOSSt6pXQpY9G8O71Xs5PsmwqwzNxTf/tmfBecznh7TWK/9
GyyTAlqdX1Bz3i3S8MUUDown4ZR90M6Wwt84DwwIJKp3LrZP98m40pviqaYyLwm+OfxveqFD5Goj
S5sxTMgH0TcZUM7YPOuav/G0J2HKzUZV6KTG9wdO9Fip/OTY170uc+EBe0DP0VUdx8nlDmjbAOla
Z0+fGDn6QJMyT+42wZXIssMbtRG4EI8A++o6GmQ1WJnrHhfib9GcF+bq3F3FO+zoWPzWxggQcWAO
DfwJZoNLPcIpVqith3Hx6DkBZPVsR5fk5ldVL2s6ZanhuWmvHLwk2Llf949s2/2HcembJzMgjbEP
PqA3SDMd3oBSeAsKiFnfFz2Hmprv4wMuj1OtPQuq3jUg1mlIAq0Hto8ic37rcsprIZ/+Qs2is9Th
a7xxqiAr3oIvF8/I9QLLnltrKWrMXdMCwIpMAKSl+ONfNECNXsalg6soWs78l5M3yN1RwPdaVb40
Qd6d3YeoV9Xw6VQHgrTXlW8yLcGSsUICmb3JHJ5vH6a7j4vx/EXgHO/qhmqyt6QG3dqjtwZp8tU6
9XdWZyaTmHLTZQV/4Ni6Mx9ItFNvNpRHbYKDHRE0jIhBCDDqwqclTs+IJyWSRqeJEdUM9z8PMBx/
kN5apUopHY2+vkhdWQwUQ3oR7XskFS1cE6eo/LjnThbrIr/TmyITRDCW1kC41a2pOeqDD5Kl6x6r
HFPARtAASY1SwAInrh75fdaXKCf0fKtgkCoEAoB1IIZttHWvHtAl0JunOJfSUBRtPlDsuotGC5sg
ShcWPHchvHXr0hhpQqoWSB/JFHDX/70vr7mXewf8Azk/qI6sF5+4Di3HedeuaEe5SeqEh2FAqYGS
aBnd1Pba3V4A0e9JTPyAwUZiGuglFdFD2x9HekmUcDVllz6huUe6rVEcc21Gh20/IqqCS3k9CZfa
JuZGMYqnXusnNNqvocPXT9wiQ8yFZwYWVVXp1nqOK+s3hveU2Xix+b3W4OLEHPVhG/9tD9X29TSI
9vr/MeGAgTSpKnEkTILHL7cLv1yrkW9kmam3JXW5vDcOoo/Ho9XIy9AklG33GCbZ/2+L7R/h15o9
OCSMIPe1wCb4LxL7xIdT1j8QfG1KQVXfcbmCDVtj8EiJaVLxomvmqpMlUqgZ7T9Yr9VDEvjmjPq7
Gkl0hI3hMmkN2hTT175zOI7zEDgeNH/Eg8fB1hieFLOLvMsY1OW+l/pHVlgI2Af+P0AYasblFa0E
KcSr2GCJoFlLDaxKWCH3ESOa5bYAVi6svU4QZ0WLVafbIuzuKuI8MluR/nEsSDlYW5qEjX1bFJJU
KdfLb9RlAKnr3H354qRhB25ZVAD+xIsaxZxD8HxMMkncK2bQHvWzLxaf8hX1/yYZvGR+1Ar5Jnnu
nwGj2FghjV5miUvHrjBKk9KGhsAIXCqefbLVahr2tW5V2xEPI11427fQn8TeLINe7O5Wc5BUfTmN
l5JilrydPGNc13aG/P4Po86mcFSs8gv/QJvsXaHtNEaM56I6zt/TTyCwpGg2U/r+f0oUAQRyXUeQ
EAynO2FkdLF86BlNCvDz6LSSRl/YYg3MNNNJs7qi2/epjr3PaXFGTaTJA+v+X//P+h32Fd4HMZJy
ecM62ploszr3vCEsGrNa+W1lBVPZ7DvRfpzXrXJnInQ6lLBZq2bSbOXts5vuQuYtW+W3H/d2DB/v
61eW2gQROQDvKcXrL9/QSu0B060dndnShfBOghuwoyXg6fUyjrnNflSHQpUsg8fIoD34Bu3TT3Nb
vrLS1z9lYYaCc7ZaHZOimYQ30S/lrIK7Ob4uJsycoVJcPXlagRabplisKlE1c6rX9P6750GSSb9p
F2+o9kt/KRMP5roOvzAs8RcvlrPpbzDX4Oke+9qytH7c75W0QnzL4ebC0d6XcUgQuPAujxynU7aS
S4XDAkSKoMWRN6ENZZLlyZ24N+/OArSKuDNUoW1w48dK1uUiDUPtyYB5989XDprc2fRCuKfhEHHD
P1HTpFBbI+7mhHPGuTc8LUN/RAVT1NpLf3kdmyUeZBwIYKbS6Q8NDMPjNyU8IQAmnKNJfyieX63C
VSV6E9z6WQrzPklSROcdbQyW5dLfvLVQDrt68kpp+lMLSoKwpTSuevXczw9Tr7FW8lq/F1R2R4K0
q/J6CZ+H2W+jjDv2h5BGPUHyXu8DFOzBpwMLd/mOffKX2Ddwr5ukqygf68bltKe3kbQ8FdP+UE2g
L6DBzS6vTmeUCo2Gy+Cipju2YOC/+TbxtvMZquT4uNpo4WZAvfa1v+kmjcbwqs85Sto07Wdshx1/
LnQKpspC3rYCeb1bJO3qtXBQBN/4We6S91B50cq/wrFF9CRgk+1xtqRf5dgXdCtzTH/EMLWaN2nO
tIw1UAP4JhzpF8pmNLfdUyntFdAv4OOKzlUCu/FvgMvhSoQQlD6swzeUL6n4AJQB5TR8BCsdoau1
KNuG32szWEVbWjUb8yGs1Qiycp+vCDbSHUmnqUHnyygXkdVXwRxsFXgnGhkFyH0wuKGzgsAQCNkS
GUiDbPpvAPnD8p0HollSvTdnkHrdGbJK54MaUjJMBPkgxJptaCTFb2AodfcGzmHE9k+1xRHKvIuF
53KV4R3nLu/SroPdwT2eR0etbrBUuCprTmU7a8RYR204roAy+BCs0LS/Z1+IdEIqhrAAvO51zP8o
PglZ42xkejm2+14v0d8CihlmFP6pp0HYx8wEoy5crPxuv4wVZxor12Dk8y/beED8pw8dXcgi2Np3
eulcE5wG/XGKLWHyMPfd13IrX34OjiSC6HPvdel/5Wsg17WOZgFXv3ZKu4xnd6P/AcUCA23bu/t1
GbijD5nN5U+u+cMnvoT0sHvbzmLlnzAww/YCD1gkLPKE0N1DzhFm5IR9gHPsYo4256vY1hAXxZdq
hskRdZBxaaG3wDxDH3D2wlVc72g5T0TY+DLIYSioqP5tTIB9SPFKFTo4JK4Od+lcHYiZ183Ix06N
lJhbUuD7hRoPLQ8KE+f+UHl293/l+oVGIzhFy/h6aAdGBoFN74tuWQm8n9ku4hFkyyrqsO1YjMwI
IoLopD2yL/ecLGjnZh97x5vRfWyNx+JfABqIQqovS9KXOi+wmqXSDAnnY9y6PhKRpKa6HhBs3Izp
A+OxtGW5u0l0U/mOmec3YAWt+dnG9IaIlSFT3lfcdfMYv80oOL9p23PEAhOjJ6k/OcKwKnW1jgUn
8x5BII+zKEnjvQkphQr5KK04E4kefoLXpYZkJVs+h9sX1Mh1QVEwvv3/Ncwl54t/QbUIsTMX9Z0A
2FAX83kzPYqSix22BrsZmr0gczOEnsFUuLZeUtgjBZ5k7517c9Aa1D/h99QDNkjpZONRbLUFpQJo
SSSgOPXp6FYQ6FYGh9rdxyX+pk5v2ZHjvyQbkwCp/9824tvjgfL6Q6ZDkmspQAZxrYffydXgFgM5
SKklJroN0KDIz8syDcDW5GH0n5MlVY33k1jr3p4NZzAwoi5zrTlAxEUzQSnnhoc8L/NcqcqpMiUV
TsCTigfcCQlib4jklcQ4ldamf99EG0rGsr9i+1HnZpGBCF8HO3aG8ZzFAtiaQ6tx0kAgUQg8C6qj
U/hVPybaQRARgYWIKnrXLlKyO6QMyRXu6mDixSYW543sby3E0ne4SJQ0x7/sxw43SNVYQTszYMqC
z7ENtgyWIdrfsS7dM0xBbrneW/+8+tusc4K8nIKV4/JWbb5jh2+6BnCoI5FgdCUhFEx3Ruj0IOD4
+/aFZ+Jhk8gfPjOXQZj7O4vB/T1IaQzIxNeyKrCsT/yw77jcykerSrA/07OLElOPC4dQ1o0Lo0qB
X5cCYVS6XMm2CQWgDxg7r84WFpUzWZy5CkdXtMQhJ6vPKGdqbCzT0SEq1Eq4xmgu8CGZhZGNpiFv
5H/QJiPzoQ4r6v0iEUNcQGXfzBc7ViKeujvudd42JyDYVmhCp64ZpAYlx8WjdtDygKz1rH2q2IwQ
AcbnlXIxoS4pADmlSUAqLst5jKhczsz+cAvWD85g7IoOG2TfiQxub7/vFxl6VKpldQw690/07/bx
KEK9RZMiT4MbusVPD46epjO/P55xa8tmE9hGZfZweBsAJbBLv44Q8JN3EBdS8UIKCTn0lcvayVeZ
lw/lzXbc7mi+QKueBR9f2shGF1HkuxYgQhNsoReBQeCHz/Kj436/iHnFUqh92tfalK1LC4F0t0Vh
b4qkXoRCYq4Bhl550FDwH5mZIvhUYzseS/MI8VYRNmYeHgi7q/jww0fxV8RxZ9NA3/DFKaGg75Q+
xmwvH+iWRNroQ5aM0TgnTrrYvOKEoulrYB5KvjLUwqwnC76kq7mIzZaqb4JhAkiaX7pTGwPzjGb9
y+xIFIonwjUORD7nQeoXbt95lRGy8OR44UHuCgRCxDf8tJdBjtELil6NlxFHTL1Z2cF9US+6pZTl
opLvwj0I+X4CGctyQtWiRmBbt7fyrh24OQJIzh/PBegAhT8g5g6wEcLwFlEr/f+w2k1ZDz1YPO2F
SAZmtS7UOC5ScTm/lbgGEwRKtcDXAa+20yrD4hMRiGm3AZYZhktHWP38UWjcTPuOGc5wiivHLvEv
52ROMPMGeS24GfIbCQ+/ypD3/BYLsQb45mKOrIuxlhQ8CW9JaiEycYi+ygQZS5KImjiWFEvOOUrh
twxZrzeLSumAslv9r63j87UGSgkFUTPBCOXtz+4wV2FKPVPRhckLE4shB2TFUHavH0Izhqerl21Z
peKh8lsFBb0u7it2z7g+sv0+hT8C9yuBVHMg6YwC9YdSeDv7OgVZyXK5cDJ1tVEpchwLOxj+JiMA
D7Dp0eUoE8vpzYI/OwNHD2JRuZroUQDIBUKif1Apvgz3dn4T/WDoGPE933HKRz7A9pU4wyVqcoAa
KtiLOnAbgYkAD/4FwmqkL4sEuditaUOYhuFQCPHrMTK/VTlBL4HU3QYlZg8Rm+EOfJ9Cmeg2aS96
62e81sFqinmW7fwAzL0vyiT17FcAsZ/u0mIZSM4YuSSVszdCokOqG9Vs+GrqxcAoPXLl81eJKBV5
qPS3dFLajbeJ95qkl5iExajWY17Yj94KgyNX/V93EWp8kP40/4NN06T3euXVFIpo9L1JB9oIJdg3
Cy6FR+rG13iuSkp41Wlg9pYnpbz2aWuv0wIeytz6bbslbVb114IFuj12hG0NQ5wHr+PECbGswIre
8FbL2zzrq6pQC03dbXfQS0ICXBvcrS87UlI5JhJDmB9gU7ZGmDBVxS5534yeiUArC8KXhMsdbwY9
0MOTiglMIhr5J9VKkWXVZ30lfhhVOihuhntLT9n6yPOpP1VkrXNoXgtL1ZLZ4o7x3Tzo6VUaseyJ
PemnwKgfq7n/YzokwaLTXOqN7J0PfwBTRgdlPJmcL0tv/ZipOrrcB5jFWKDBVkwJ1/+JTe0nXAt2
t1lgtZ8U4Bl+BSfPfkuOsELoUyw1s28unVyjBnPJhE8bWVGYOUdD3WdtOqMHdXjLKotlwVTRvqEQ
evCm+HQZ5NR0R1sI8eaiawma7sPu8WkYplyyhJbyqZShNxmKqn2ZjcjDNFTWhrfmKpaBSKPG5g/z
osgVTEwM7kHLmVpHuh+JZ38uhgoTfXQHY60TS8Yy5ai/vTmrSI36puVDWxNbAl1rpjDopAx4U6ix
g9msuxGRgK1ocNtL/YZOPjR0pPj6oHdNnZnxTWhqw7lc/EmHCtZWNlh/hv7kAs3SkhzDfNCxWNUi
HUfvsRnhUpf8FGnRD+qxrTfKwSsq9iMl8S4gUM9gaLGTJBXvFYbvbO4jcraxrssYTq48micHEdlo
OE3u/qbfLgbaW7zd43n0p5z1qw62wVY2UHhN63abrD86dl72twkpYHCrtmjH4UvaejqWERgOAKGs
1x1a3WRaGjF94J/uJtO7XfmjASPpnMa+hQK9/hP0JhWIFn/ABj5X6sMk13U7VjGVy3wS1wIDpGfj
/lG6XCgLFguP55K2o66C7deUbkpfbDi7NGSwQAyA2a3fPDFn7tTxKgXDXiRfI76N5jU/bTVdvVL3
WCRPW8/3nGfvJ+ENB2mTEdq6sd0xjFLulKGHUxMYGygBxVdo+46hSrDiWf2iy6pY3TPY4n78jQxt
1n/nO/JleGWSCtXKKOtntcs+MUoMfymkwIkvMKSxKTRIWSpBISFCyqEu8DbnJIuQNuo84qi9iPSL
sLXPW3hroYgET0xlMcrctMjAzFgmwC0+imQm2dMyE6mV8ee0IaK60O9cWpf64sDM0lGkBS0/ffor
fZ+PdtyDeGZkzliuH9VweEYOGLn/K4iscWil4zRYaUshwwCueXl50ibJqpmFDnYLUuYcEsfMqey0
wBAOabz8J9LcKi1XAZfaWjxJkZ6Ii+uhudiGidFHRpALrwr3cD6DcQLdl6UMVZ76IuJmdJjD4aF7
XVXv7w84bcNMEmYy3majChLF6Ml2aXt4cysr01d1Fcow3r1i8f/QOjUUmEy5RMvNFBHXXVcH42ww
B9hQuRMOZFzjvLfXQA3rdM+kBe86y+sbaC6aK/mX3apszcZ5YTvfx7cLsf2t5CJ3GFfPC8fxUNaQ
R/gnMKtNExW+oEXodE1D+hVymDHbUiGHS4iHmnxzYyoh2K0GNcIhQ8rd3vrVi5F/rlttBArQXMwz
WJs2GPdzigSjbM9KRSt+onHeede/IIUKNljZvS5blU0s3e4am4SCB7PRIk53JkQqGhYXYpuxK9ob
5UmJbmAV6FuPAtBoWMdfo/MNqJXOS+PW22mQ1SxwofrKzgp8hWifKKc3D+mB9DuZa6C1qGMSDvRR
w85Jfi/wHKY3u36XNZ1khyzRPYD1KZ1zttYrQhYPqt3W5PDF1qSX2nAmBHEkgnG2DL51AlNsnU2G
ML+343Po3ypTGyWEYQvFqyYEBOlOePJuY90zFRdTTZkTLiHJMKVn6wg992PqI3KEvAxFo4Sq26gO
6rJ77Ngcp53PXN8Dte7rq+UmqW75cGep5GS7j67OKlVUmTZapCEpSGJFtMxy95B4w6FDF9Kcg3q4
1FzW4ijN+oIyLeO0POPSmEh+je1WDMn/x4w5qlcL4GJPu4IJoYUmht/Aj+A7KjJAaGpeSg8V79Bb
iAIcg7tUSY5dkK9qrtbG55vhjGZVUyS553TM7zT+K5VpysDygPYCktrEeIsBcNGudHePTxQoesCp
Y089jCNQohSKF7xLJnJkLn1RXv2pGKE3zgU7YRPGw2yxcAL86t+r82Rl+KibJsxh3zLRWdCYaGv4
xCXx9xeUs8/fjRKDOzVlSfKkEKLCQTTths52ctnXzzXuGq9hWYy9ufcDh45Tz+eZC7+mpOqljWks
rego0DzRmPZg/0l/4+ML8xDzRGcznrlM9k/O+edJGUF+sAo0B5K4dH/rN8CVIJY4qgOvG2S7AFO2
+8dwRyqJxGbxrSd0gwlT0LE7l1qgKEMKm8qWyzPeNM0YOw8Qs17irT6BBw86S/4se95t3zNIobBl
gh5URPDbiNJ4sEZmVKrXHfS+4vkcukltdguFwAQfSoIoihZ2CQ6Jkcniju7kBTckZE74h6zYIIcH
UCoQC4enYpnuVniTDPa/BvGwTpY99QmI0yY3oe7+JOsVHUgv0oIhMI3XIY+zMtZEprCDMt40/7To
7dvST9LSUoVkHZMt+foGcmfNxJNmw+mlFdS7ttXOauZyS3ZhbZV3eDMQOppoYt1h3HirXnj1o/mu
tiJ1o51JWroZ9aYAa3BuekMR6fvYK1IAFJA6AfEKxwZ1UlFJ2ae2sGey8GqvzxDdzuhgrYB/2KP5
km6wZIXVT+vhc2hhWTgG46cIe3W2Ei0z/LQn8JEuolnhFLsHvYu6XEPJKTUOd57d9hguUTdT3BQr
hma9e4AePDeACNSjoxQlSGAUmT8hWLQX+T3dru/fDoOeOIs3NbE+uzLtewe5KeNajuANOVwqFBjy
3l35M/ZgKp6RuIhEWaund1DPEuGc7nW5cwc1FsRopqbmVqaFJZECxUNdySGZnRjWblXJIEdkIOnY
M8+/VEtv7uWdwueXUik95YJDguwzHpt62gVQ3VdBCkUKb2XJOj4MWtdom9375WQCLhQscL/7XxAY
zfNC6hGNPo9SGPhWW6UDcskPOl4Lsr2wNrKzIgUvwcu3r1OgDXNOzV1R4ll0YMr/Tj8Epgb4UL0i
cE7JYk++17vKo7PMgclMtR/cda3beFrB6IQ0sQsiuaIJY3BMPRtVOqcM8sxsftc8w3p8NwLzcraN
ACOc1CZC6d45GFDCJWBNZ7D6AboKyJV2T1osZYNfTcVL2jciRsBgPFhxAIZuorbGsEVW5HZZ3axx
vToEhEIRGP8n7RoMeYhSwepdeUlDDC3ygtHk1JEfdMP+0vMZtq2sJzIa2ADm/Ceeh3LLWl8nnkxp
/0/dYboxsGeGJJTWMGgb+Q7XYIWqRF8/VFliB/48VfTmoGY+Zre1u6znUKlYZri7dkyb3iFFVxi3
9SMFlPKW0Paz2//XZr0XWrrAl0vCPQgby56PRzpu44vwzpKoJNLwlWglExp1V8sgZPacQw8fzMta
DxMIhdfnHy6kXpdUftCMtCBeEH7/kraPNh4By5B+sO+ryI4Qrw/A2DdZCbbgTTSLnVqxudpATq0m
pSJMvxvE+NRQGT3I/tmL9A+/eutrrlNQThvPeSeSu4ifDUM+n1CjwFYswK/2bao4Kz4iSRMDMNQN
49BrBSt8r/gEXBeYxdM6jUQeTkGvFUXIA3q2Sj0hGgPjFeAwFCYjUU4Hdcrpv4MxXQGBXiEZuEY9
S2PvSXyRt2sRwz4ZBUSD6O+9C1wPv76tyBbUm7nDmP6T0a0dY9DcnmmmQPi3ZhP7xi6ld0J6b/kE
eXPA6H/BJaIfxCA8wc32F71VQzpEy+GEo95d52sWhP429ZA36mVmhuq/MGGYToFq7zKQXF/S7OHS
Ro6dEI/Y7y5/pyR6Tsv5A0Q+MNo9QcP+JBm9+4zW8R5KNxgiQy698+kwEmevWeyJ/626ea3phit2
hftsf7iYqhbvEgGuEMufLZXNMWHUIqiXL6IGvXGEPQYq1KPcVy4CaAaftv+LSp9UlTi4bmF49Ixd
6ymj919/sSe9xORk5PRY8Gg417vmTE+R3F0EeGSM1o+cG/IuRScIRyCXR86VIidEj9GqCusVDsw5
cCoembyfLblM7JqpEWr3sLrpETt8A5TBWBH2zBNxPdLRuzJYULbciUVxASuIehDuHw6tDmrpWfrd
i4bf1+Foe+oQ9NggmvYUQhN59V4U7T23w9G7xmjolrIImSG/5XDNFli7z7O+6976p5ynZFgELS9R
N0OP52Jg7m2mXMWkH/eWj3t1zn8syzrAZbB9qJOX+4Mhrz5YuWu+HfFxC+EjqIczxgfjXYCgxLsM
6jgAx2KLHTHJnsgPSgjl7ZNocAAJ2Rvek7rSJQddDMU8pi/BDLjxxDTQrDJ8uYxGvrDqLhIb7UV9
Z6SEtXDusSJRkDsny2oVDsvYPSvRPZFcQ4pSBT88Q2TUhpptfOoto5is8/HGHZNSwnwlj55DCQqA
7ZvzDiPrVeifNI2JjDCLcGeH67wHRKHHjUBrMDAy7S/trDtVU2ZWMRfzXgWQEoUIyJrnB/6OblZD
BEkqa5fT5Q73zSFvuL+kQFQNxko+N0/2NOnKpTWfgjB+aon/GmHnioL9GR4oresjopSWOrO0QoN9
LyL14dFjHh5gh4nrutA01uFguUUbB+JyXeqMkX733nSG6sfSZ3btlNso3FGuRLj8UDMt2a/WBCKM
2AlGvfWsOtms9fR7RYNc9B4DnR0NZp8yjR70coRnvgXrPGZoqQKRIJeMf/JbHJ6ewFMdf+VRs+jF
61dNpQvXXhZo5xB2k/4l3SCIL/6YS/vC0xB71HeCFtR1obiL+Y7LDxOjLSzDKB6vPuSRU67NZtE6
LAqB2SfAt9q81zsNnH/wMLNDFjka3iV5Y/Xn8FRVZxic51hcyoQwzoIroBmiF4qJGZGul6TT294F
s8YphMW4XZVIbdiZdDDNDZuTtpwmpBaZe3JL92n8P8KJac5HfX22XxEyIHijAisSwtCJmW4Z7Egv
sXv38sDGvH64Vty4/n7Vufz7uI+6xMpMA+ZU2T/ZOGB6eq0Eq6srSjnBc2O5vRdoWBftNjSoeWQ8
HsEojb/fms6+qjWCc39kI7ePv+X+ZNXUmPsNyQIEpp3rvic01NFng+EvcSHkdSAgDWcM/4E2kSiv
JVSMRb5/Iv8efniKLO4A+Jibx3xzms2srOVUe2Usd4rseseo9ifenGJ1G8eW7G6RKTaFygjdJSbq
ZPlwObu7tWIemkf6Egi5JsJPmmlVeftyGfvcvSofTL9qS3PBaZ8ZMFt5uFir0dna3X8VcdDlTfm5
aGYmPIFZPS6cO4HGlCi2lrm+ld4H9vBTrYtSyQlXq4daZI1TWKT7ewSB3VcCNk2C1O92VoMcSTuy
rJUcD/PHm7sHERnJM7OWm2PpkwsB6xemKcWp9w5s3OVr/1nG6g1qwTmbUNTbNpyUGoWN3WOtZH7Y
ryG64dBd7V8gWpAehWOV+1NuXYyknPLSkiSIQajeBxJ75lJh6Fme1ARG6Z2sq6VE2x5F/+KCowAc
p/C5bctJN7RNBPbvVCBXpK9wVKZtLQ5lMJrCHkbMseLmkZlmpkIOYvwHaEsRkc2AlaCojx34R3JC
RV+Yop4EyzNAFQYdMoVVAQBfyP8UABNlhwSVGuzekZFSadbUNBbmQH7q8x2ajmEGtxqzHMhImLo/
0IpgnxNU4zeA09CmyADOsEV/EBjJJYPbzcpFdT/mC8b6xLRhXx53Uz0C/+39SUp1ny/62AZ3Fi9H
GVrWmoN22ooA+IBv/UXOdQZ0fyLaJku3BotslzvYtSRzsIOYgBSJ37AjJNgujZNlAgXZAUKS1VW+
7Y0FDxp8zljbdT7cPdMYIGO6Gye7l4IadlxbQrB652vwCyzc0R0i5U/xwbWpz+N/CK07o8KI1cww
4xKFNVf9FHygbrgPrd3Bq9vGEmvSjUppEqlUuVb6RzCXGXVb5QAcNllNdUYazFlPbEIEuWVNYBVO
dNJaH4Glc6jIcv0LX0tsBnM61n07m96JYRsLlzeXlGlBYRnWtnqPd+Yjw/M8jHnj866P0/jDUPtU
rvJMgwwHAVy8r33Ot6Pp9hkd8ZxG4IZKJy2gluXPgcHiuG8caUMGGiwY2lbmSui59azku2XtCC5k
2XwRcnBkuvIvC83ebRBt1AzTDq3rqUKVRrfBIBAPDgVUmlaxLESWX9sGcIM9/SrSinp5XxtiZkWg
nvZQT1xxKWyr0aG4WlweUgj7SS8j3wlZcXymNPXpfaXPloQCdR9wV54+XaT5leOgsJiVjKOg6txC
FFNSI1gT/IezHsJTu6xSpt2UaB/rgLLqW63LH13yIc20SrtZ7eP65xNW5M06SlcXNZFRrCyXbnLh
v/s0yJF0DCr67GPYjSNnEQSdOSLweU/tVeFC3x+k0QJ5ot5bUziY3pgPnaVl9yvDoPpstI9+F1qV
iotfEaVSxlohs11H06LUDizj5vDif4fTxc8kGmhERW84kmCOOKSbvAdKPwjc6lu9vuYJsESGTTQi
0OX5yuSbnTdAAqsv/vmoDG4b83zPAhJWviDiHqWWNf+Bh1Ig/Y0D7kvWez6OQmlzLPOLtLMG7ReS
a29tb7rnuWSDePSOKJTw0TI4gQf64VioYgE090uojGoWgjuFTUw/vWGtPrQlC9FiaF8YgCTb2RXq
XOZG9fb5efYJpdrk0PGtTH2E2yqmvKPPTUFKECoc/y8TvV3TsaehexAtFWpaMc0be5McyoMJ57JZ
9xCEIXDPX3YsLdvYl8YqNj62W8TWTn+DbwHVOScdf95BgVOUygrDwWOdocifptLn2XXeWZEyLfoy
TXkjr1/8WBIZMi1vC3eJcA45SgGRhpl7Bhf8Oy20vcR1KKIabKIiFEid3GqdwYh1iB+VBhe/YoNy
Pm/8zXtWOEXn05fa8A5GEe0k8J4JrJqnW38oidPmlGiH4Gt1XiZjuidjM2MjAGNlvIwl1628mdzg
1nv81pGG6e50vDhg+3xv95uhxHlM79oI7zN5aMWwY/MYvnWibddKEugtTo75Ol6l8lrvSc45jD1o
6WMJ3TK/84c9jjw3GxmIcNgHcs2coj4mBrETlbPwuiHS55xprynq7lgtXZ1tTxtpVvt1NwHGQQh8
a+zbCtWSKShO3//nZBWZusTEsrjAi5IuZm8SyprZQ2XoI1mO+1dpsIVMkHj1AEs4blL3DFN2xzxV
0dJbtxI440t+R2tFP1g+LJiDSRJPlDgMZZSofwJ0psQPqgfCEdHjdAKHTvJVf+BotHDu8TqkLvKd
0O+BAyrmJ80zWnmE8Yjl2tDGzmZvgLaKQIvgFOX8JiFLEVfTdt39cogSJdVNzo99JzbipbsbM0/f
mp2dLkauwIAUrrVNNz1ga9DCy7y9JWHm7+TiI8JeqccNBZ2Yk80WLOdZGOQjZJuVS1nNs/HzYS/O
B0vEhrBAtdNbczbaIxMgHj5prXI4SfMwTXkqbW5lY5VqGCsezu1D3r+jFxLOz4ByZARYzK2978WO
axm32FKlWT+oLiHxSWKDN0GLkYqd1OemD1PeXjck6VFMeWo6b5AwZB6xHkiXMZuAsFIf/rCpuYUg
NfShbecJGY34zoZCK/GdG1YIN6G/7wcsneDNOgYrKCh09SzAL6qYpoUma5KPDsA9Wpqxcu3M4Vw0
oYRCDHsfXaxq4zn4k++ZLFVV4Gbkalm7jnpgLdv4lil8T2WCPuE8X1NTTovCKPx6HpbBWj/NaHRA
0nGrn2RQvB/PGYHzN+lTY0EmyPa1IOugs3CrBZt4o5tQGanWPPgXZTnuW8mj6md4wVVY00+YxVu9
TXQwiknQ5XIJboWbxHt74loeGBKNYgHt9Pm1i+2YAfW5OmcrLDoK4yJfXALlrGr1qC5gjXawaFC5
Zdrg5qZNXSx3f2QPzTe+506Z9LVVHviWZfWfXTE13quwNGdYisnLF9EJAaKryMAd1qmVQeWMFerh
SE3StP7ObVesa9ermuLIrR33fKGISQ5SbogAurL/EYLA4jDz5mDMfVwzBIS3zrZfZ/x0TXYVD/fk
L9h5MAm4gVgWVrlEdnrlmBl/YC6d3sVkvVKqnnLIWcOPDNeRl8JwU4tUqTiC2EGFtLf1oEZSpuxX
cgzb39idvi6bs+I9hu89NcUe0AbL66TKw9xrYN8He9G0er+ihblWUC+OXrbgVhVzrx7VX8th3sR4
3Trf8l4UYIe3H/gbhMbhnoSmKqeiWloLkU7tUwS4XBiDYnrGJ0+4ShsxX1izL/Fm5zsFEvtQvwFW
hEWXBO8x+vbgqIY3m2t7dmPrZaLZFaOACadt0fZmFoLN1OTfh275o5amXn+orQRUCrvBT7SfeMUV
lKHqxvkOKDKKjisxH4mlVKa2XorAPppeYP/niLIOZaYzHSlUkWVFAuIkI/IWT5Ixf5gBCHniOeWv
7FHLz0r4kP9ryvpeIK8KUiX7SzhRhF9VCVYx3wMVfu9oZ3dg0pQ4447fybeIFPIbROJG6Ym15T7T
VxwN0f27wHguz4WlmARzPQPk0BVnk8lRzyGWNKSMok+pOHv3ug0vcw7Qotw2w3T7PBMREXX47FTS
RTA41+K9+6qBH0owR2Cr7tHoMgBw1sd9YZ4lqJZPStdy20XS0QqG/DkS7U8ZuWHEn7Tp+UgdecvW
Icx4J9ZrXlA84umJMKu3/+Lt83rxU/CPdvB1Y/7gFBSOm3i+dDrt0Nzqyi4GqsI7hsLcGMzCZKUs
tmrSTF8NAiTGC5+TrJttA9sduGKmH91eEvE1QwHkGptsCzS4uotGoMAdosXzniQVsEsJpgFHRn9Y
C7ea7yCq72B97oPEBzDQBt7p1ntV6OqXnzIlCKaF+8Psq5LLioNGUiYF1YLk3YcDmp9c25KM6Stw
AwefZgah1Wmln+WxlbEYewEUpJZMBUrHLyjBYHdZ6Uhm5OOoX1/EAGUlu/KwdgkyjTnWH29kQ3da
Vln9hWSqYeY1Sy4eG66qztgfWRN1rGhWEM3GGn0QQfUqjnQtdkVDvu9akVClfrMAmsNinw6RF09t
h2O9kjqpvIrbmg3qycWjM5O/jfjgkqA0HGCZijRS7oa74dAABIE8u/oS52AK57f4z/iVjFiEtXFc
hsfvVLRpgIY751cEHplql52EiDBJrObpwc7a5UG06qTrnmR1pg3BVSFXu72/5/yj7SBeBwnwUat1
MoJr63y29Lj40zUL7Ak2ItM15xAK2MDCjigWA9sUwmD0gC12uG+hiYc/3lKsy2wOTJHOkUSI9RpD
MRlFgqVfXFD509tZA4gTFWvzzY0xaoO8N4RBHznrWEtKzltwVrS1yHmlh0XR9oGbKZ+KkJaHqmTQ
DZtY/PUgsh5vCW00a6jjpfe6SMAPD5ZVfVbX/3u42ig2X/7rEkd3pvPsUP+cRqF+377Iff5JgVju
8MY7af8eqlX6bOdF9t6Kn0AATgdT/wb7hwj/0l0eOAhk3W+6177WqeJoZ8qVtIex3SYCCW4pfFeC
6E4rl9deEoNgSVm1osasb5bndKLvrfbbSN7Oqtdn6iyDvG8YxcZdu++ubYUjtQ/Db3boqXgrA4nF
JGQH7T4tXOqXCTGBvaDM6ManOUffxpRACHbqRTHDSf2vWo+m9R09HikeZd4UwbKfjgL3sifNRYH9
dRgFJTBwUv48oVvwNooffUwrpBAMJj6GW2bPL8e3fZqR7/ZQGEfLW24Ga+J9WzOU4zAJeRykTUB8
eUiSTKyqqc6Zu1OYkrGK9jRz5YIH+VZ4hyPfl8lQWh7Mmd/DFUuoqMuubNY8BmBKpxEJbi1etLNB
vjbeLzcQxyIetFEGFs13XSBBND+dU4U0Wj1V5DCzj9bMKSGS009GH/vra+k3JHFc7YzDql9BsKBG
S2Lfk19R6xa5rT6FELZqV8pzeciLwJ6DHGEazA6k06gFCIxoyTLS/eXONDLdHIJ87B2TBeaKPcjY
n7YC2Dc/VKaycFk7mXQeGOyVKtJrMyPUHH5Kj5a2Gr/YJLSylPZf4UtXfXkmI8S7eCFtdYe8qWK0
aCMgv3kR0jlDKCIKIHTDFcPbF73uWLx71/LCXUDuxxfsBiBrMZDqS01iYDLEVUSDe2Ha6JVayKlW
NNoCsQslIZh+pIj8LcpXUOKLdXwDuYhsOzjbgY5HYe3tYF9RTc44gNFV0paX7onpCJbQL7An34k4
bMUUCMouYVyalzjgqSLgTkqz86egLgYb0kWz2h5zQQYdLTzlYjrwpyFf+Ko2rKm4Q9YtvybQOHc4
46VXWLrwWAWjz53+AInfJta49pXpUe4tdqTY+63dIpTaf1CoZA5cdZ31eioJaTSEkYEZ0Tt+F+6K
Q8uAzP591D7JmCkeejUDGzVhUe6Mt2ffJaq2AXlv0bcjgqV8fedRNBaKccRCcAawa068km3qJTt7
5eSCI4bu1QByiSWMoW6TiM7dsqHVxJNJ/dUIkSnTQ9mL0UY2+TCnWx1VSjHA+6sXhPNuxzT4Xz8L
+inF0rJx6EBkLsmWYtcJBe6QdlkfvdxOeIeUxigb/LaRjiYTqAhzZjUSa/BDRizz7hdg1OcuzYFx
CrciMM+JjEbq8IkRs5wrGr/QzhtqPYOmKJYx8CSGWveiRNXIuoOfSt90LUE/+p8jpJ+L9ITR8e+y
69vv1ku0ec4uwHoZEQD7i3g2XA/Gda4dcxt8oRjF7WfuZDx5eRxGpSpczcB/kyrycVQ5SjtYagr0
BtWIUIqoYKobPRKeBti/S/2XsApddMMC/wUvvqb6VEaQzoOXwxMUfTs+WIS+rll2oSdLjk6zFmW3
1tG03AN7U/jik1O2K6dPcx5ckeqaGAXLMqS9tHwxTwBvz9xqavGqvrqrqYWbzbWnqhFtEDjY0chg
fGDBYFFAuxawnQpYzj5CGbeT/vbwNX4xM5afzSNisPjjZGdWqxSkjB9wz00WIHL4T0ojjqlYD4hl
9GcWNZQacit3410fdNpsVdk0p3KB5Zc1nQmkg39BsFtrvods67ko9tnTGCeXtIbtzTQ0hj3KdV8/
UxaVxR/RIBHIat8+iuuDc1dqk6nF96fdqz+z64e28DdtbPOEBLpooK7QlPWCCUJJq+HaZ/sQwIVn
gWsJEvRim14QzJJoHjto0TdgTNcpyNr0jwspDGesMNb09xjqnjyZ/ElFBwhtWXRut6DjLcZSkoIf
U//liQZ/FO/A12oJwNyYRzani8QscQumRGJ5sW1lQ9jujNVOAnAlMFdorLVorBXtyWo24MoVLcln
r2KSlJQ4m6oa1VzQWIA9MFvJ6qrMQBiNEXhTTQEyxWn6xMgCRi8LrkZMxZ7N0D05d3hQ1ue2o7iL
geHcYJccNAzdOUp+YoQ3JKU1A4P0bbtlfEd/lUIAz2/n3zFtIWMHb+eENxtiUY2uZdmHRyKZWjZN
AcNG2LxY7hf7SD+hqfHcRZotoi4cJV+lBT8eWPBDRWfFzRjNqdFfCX7xLrZXCfqQo6ivDdD4Homu
GSApj0ItIzjMy4XLv/SDorBkFc+Yu086z26TpvIujUCKtXC/sPwyAyIktINgoc1pVNUpNqjCpjow
qMjC3oMPVpzU5LjV88agDX/eZF8/8P4TU632jqWGrEVFJeV3RrZEQ/8uXsmaglrfaEm7zuQLXo8c
YxrDFncL2FQG0ezDYlAaDeVmGhJiKKySfYJV8yVg6HPPJszSARsL2IKyEK7u6NF8i5Vd1WY9AfOw
YqYhQr3QTOESjFtoa2FcKPwFxVnYNCZDAqE516xCnM+tvSGYS8uKz1uXuJb/W8foyeRQXCUa4xp1
fmsc9T3ehMjm46ZszZTn3PXJgVLMcso/sG/v2WIs2CWlNejpMKU8lXfNiaiaiG4UoFSIjhVendI1
9Bd+iLCotjtz5q453eYJ3XTmSVt9/UQbvaCF4qpb3Pj4gP9q2m2wF9DeuYouVOkk550dLnjOEtqx
rSrCKt6LFR+r4sTw654EngyxuLcx6B0+xJqL6y2NltnzOZfz/eYdcKOdem4WPVfewJikyFZKa2tI
lgif+LtIskA/ttEg7wumeyG4YAMlOvPBsUSkP3TMhzfKYxXeRvcgrVo0dg3aB9DOR5vxHVxUL1P4
KaEPVRzC9olzsb/2hgJ98o6W6ON/ZYsBaq9HRcupTrQcxKaNxeRUFbXSyC1wwvTjQGEWemY0hc20
hyf0Z0/HSNXZzd4aNb2iDqbSmZkDiJLxbtjeSvCJoMBYwKYd94Jrff13cnAyy+Y3GQGQ3/guay/t
XexxBCagW6CW2BObtAXIKRjtQr3sh2TLw4+vDCwZOAAOq1jOpEKE6YioaffHyldNBSM+nlJgAOdJ
dDPozGo/b63f6OilIWUKPPA9bcMrPrqxiCi0m3A/qw+YlVpGCEBfmOWszaQK7Nq0keJuVwDQADkH
AizeTpPZa1195MHl4YxdtFEQDHHO2dO96zHs+KhknAEiOLoeEEeefe45x9pm/3rVth8+VrckbQHh
H0+Pn7SwUx4Hl7pYN/eJiUVi+UBdrajcflOZ3vuxzhZs66KeRnP74CfGm7CUACGw90hy3m7eUxjl
iHBIwHnxVA4LMghh3b776JLqbTPjXFAaBS5qBvNhdszjnOaA+2v1Amy3bOYPCSIjMoCns+wgjB4W
vsRosQo7ZL9Ky5ndxJtmo7zMAQYMKFrdQnhHR8niKyT5sIf4+qDbMLOfTgsbxlTOX2Iv/VMsLqRm
zw8EChVZX0td8AjCcfI6YYILLOxZR0e+ztEgSVdjWF7zxQtcvJg9JmJTOpgEcML+hiYkFFvtbOr+
g/RxtCEsh6eyCxo2VSeGG+8amSp9PFvVIg54eih2ISP2CFRBdQj4MwOq/ZBfFw0fCzznjiHWQyX/
aP6WFnslRQVZKdyJtPZcAuT2Ymkrr625++mPb1k5rD5D0R1MKa6AsXs4ibhxK9K4Dc+MJin2tHBc
vEC1PENOziwccBppmdVS1IgsSSvxnmB2KlXLvygibdPXFDplPw4YNQc7X/yKrtigJ2PWMiywEm+K
3hkNmsuQfTQHHuaUusQylvaoSLUqajuNFnakHi2pnuLpmbfpD5QEZJiGmJ86ZT8Bjo1NsufDmprm
32JwN9mzynQaoUGScIVimGRc5wCNzngvDl/l4tswn6d+2aQtodUjtrVQdwXhomhGzfaj+/sIYmby
KSYSNOYCQ5TLEyAcR8hNSJxMwiRN1lz9bvFXSrwrazKyMDOIHoroWTe7OWCuAPXxUNiYxCKhpKM8
va7aHsZWJ/j2R1tpFieZrRE5KNxu0IzjHChvZuI8d5E2nvr+8EgH8/4VvxLXVQ2R5UC4OYgM5d7d
UuaOQikT3p6djHluv5P/Yg9QuRT5nZwgj0VSAZarqq4KhYGc+jZCATmo2GDMhce/JJCLFa+la4Uo
gqXOAHOm/11ISpX4cMJsZ5+Bl9q6/Cu7Ix0XzWCKNo5msCyBbKrzKXWthmpJzxI3cNuyznD0xaCN
2z+4jNkws4pzO9zH9TSxEEG5zzoLQ4FNUJxpZ1LriRnGOExXdSeDLQEJfMaGpknXMzOgqCQ4gIlr
f/yHQOvTlT29ieccexBqayL3tLCNTH2BobTNX5Lb9lwj240qFPozNgdJAXcOrzs9Fp8l0L7f2us9
zkwtq2NDfRe48wfzRs1KssfVc8IFxVVDDVecy93TICn24MlssWvkMvCYtqTtrkJCb3JUEUn7TGS6
PypErmLrW1zJ+eHQ9rZPIgfLA09vPt2NdSF6yd8xAxESyQfmBad1yTuqK+WNd36byEro5JGfrzGS
h0zeSKlE0sJq8w33cOA7XCLi2u5By41zllhK4cXxX5ef/Vc2SXlo47/qZTrNt+xEDsuRnDmi2Ka+
Rl8E68aZrGESKSZnGI2PY+Gbrra5qjVaOJ5jZPsGErNOeTzriM7iAyEjBanfezLkFAUIZfAQFzcA
nJAvSAimX0WOuzIRIESpYLUgVe52WZMgas4PqBl1w63Xh7ISCTXFblQ4tUl75E/DSmQ16cD/PvBI
khwSKxhHsluQQhsQ14IbHAAOhRFeQ5/Pk3d2uwb+E9i76qV1De4oK880WSMaKjy2Cvgd/uODOaSW
gwbQ8rJ9UTImt6BatgvbCqqSHZxOlYaD9ZcKcMlf/CP7gsjqyBeSIiN505BEtc7wQNWCtoOXslXE
tRbkkZy2doCMVxchyc1ArbTQDGrOV2dSkvUGxcV91mBAFSEri+EDXgfEMZZUx+b9zPmuDoLgjol0
HaufBZdxZXUfgY/GQaRECGhEticGC8ZTQMuaSn5TmmqEo/mBazm/FsSCjYAC8M8Wh7zBKt5R1mai
rYo5ckIla8+qpjfroqz+K7QOTBbMdsQ2THtsc90RNC+bEfYnnwYW1qVMm1wyAq+KuCPI2S5I7dt3
xCC+G72OphvDQNgMy3hccna00+s5NJsUbTdlG4ISFPoi3l2ygVahvqw437oD2hX4PrT4FlMTIn/4
W/EVuiVTSleYtsJ5SPQ9ajrlREjTdrhAjV3/TGLsjhcgkx/MYwY9VO0wXuuUnLDcFQndhAJxIgNJ
vVaHnqqtANQLL5N5c6IER2Hlf59ByKH0mdqE6AgRdT1VBLB1Yk0UnPdUAm29oM2KWiGzMItH9Vbv
HSKjy9QiQVOmDKYWcLP4b0wUW8yeYism8wC8NPiNTpbszYVLocw+UJg/zOaB6kqzeMtoSZ+Mfiu+
d9Or+C81RN3/TUyIwaK4x3l1ixRb1lCp8dmOkHfYr/3CF6oUkRUjmGg7hX0orY2tYVE21RpXgWOW
8AC2M8kQJxcN/o0KnoKEuQIN2jBBjXB/uEgTPMKvzBUt7kdNESCl3c7vuTdjrzVuh3XBaF19Us6H
qq1wDG+PmOfumEqPbF/LJhh7q05/rYJTwnQ3QgjrD6D9AazSiE+mcExz8iSZyJamMznT2fRN2ohs
FrYVR9tJuI0Hqj1zn1qg89wvPusxhk0y6I14oeKYU3DV05n9yjQtBIPw93u3rvhu6YeqhVeotaLz
NdC696t6+Rn5On12oulaWZwpxPTc2IgFN/OPDkmArEumZ+z2L3gssnKDJWlKvyVCguDUqSQIvFJX
UoU8hlC9BI+XCi040qLfXfTmPiDUH3c4iAnHahr1337bEIBFGaGkRvj5wt2lqxUJdjUOq5XBYW1Y
DUhupv+JDuUyXgy92CBqcj9LYnU2e4uytnnmcPbIL1vLO7KNSS68G/2A+FY8DPBcS2adl5B1PHtT
6ABHsh9nIXsNPa5aPyHwMAplwFCjSruZNxmkLRhjiH0bEI8qYpFk2TREu2VDFtyp3a1mf6ySr0GS
UJL1NlXv00sNz+XBHvx23lmVXjI2H4Z1uNW30oUm/FxloFZutpVLQZaROCjfdsABXhp2UBcQcO9c
1RIk0YpaZ7JC3Z4MeyP2OVRTsiBnAvuW1iHECRbRy6n/OKWFD/wTa4/Ww3bH6/RykVo16iNk6W77
qT+IE7OWdhPdQRn4raAoKV0uhlXgIKcWdbq0cvmwO4sxAzToP71VSsy4Snfo/w2XzcfNUNTMR9sD
Q1FmAJd1ah2Dz7bV34psMAkNFJ2A9yQEitzzcEhX4v1B8Y3UvcqNhRcJoEZG1aQxzkxbdUUVtGe0
OYszK3A3p2jZrzWE/37Plys8xOCwBMgDNLc05g7XRlDN1a6J8tHWWyfmFmU6E+H70Xb7OVuUw/xr
m+K5g04bT6+H03UZm+WRL6r3SXzQuBI0c6O1+sZxxRtoKohbm1ixfQtfVQvcY2aaHaFN6V+tXPJ/
1deDz4J/fr4QqVW02YKFpxtaQTR2ZY/MEPJQ2zcSoGELOqfXiz6TJi+0dmpoRdeAw+f+JSuAKk1/
8KKRsEgycbSZexlcBTwH58c3y9sTd9oi66k/F7kWIRKMf70UFbXSpuiPtC/qCGSfB/MuHlap1Z8w
CMtQNpdsh+yokqaeQSAtwqOgaNS71tgpyucl/+nH6y/BQuk2M/9uGwz2DGDq3AGSQwdf1RM5LXSc
5d6+Pa9+73DLp2ShD4C2XkOgdD7lnXCR+7cdhvFndKQV0CB73E0OYt0CT0e9JONV5H4LfkLnE4cB
2OJ2A6waRzDYaShLJQqUp3AQv7X/QLiiULyywtHT6PtV0kCc+9gU2pdtl3W07arJqMJIc+xkmfHD
C+2T9ltxgxj6NVu1R44pHMt/X3/G1HTBJHxZdWOH1DMaEJ1aCCiMSjMukKbggiekpkIcnH2LJnyS
AYAua/xcIMXM7U26h8bNlFrrV05NUTcYCrYx75kgQGY+72GiuQGzO8k3brkiePGS+c+szRLNbVqR
Zisu0VGrIvxU9OI/oKYQZo1BgxrGrQxcTK34qGK3eT1fz/CvGfwRzMIug+93VC4RqAazYMiNYoZh
qwPy443l/v7sn+yjnC4VqbQGQhGqnCqqj4qKw6igu9V8OQMXagiuHRAsES9rJLfw+Cawp7nb/t+h
eCkjW87GVodOSkMb2xRjODCBeHiX7y0pfTbYcRD2VDDhAIDUtjGfBkiQHw45OxxBZSVVWPcW+lp6
A/VTw5LE+R7Xj80aCw3KyYme8y/71Zp2e6RO9pjII9ZvoFurxU95bOCjaI8vL1q9618wPEY38v8D
xerzGosid/kM5FFoTX9k0dSYDNM5huDQzURecdBqTEyMtsUX569qqYtn/rlNj7vmUZ0d+hMr6Wg5
4vp8O8eEMxlc9zf63DNyzG4lCqcUAjgjkbBfvX+Aam44dFMfn2dJpeP8iOTFt11EsLj1oNKHR7JA
B9f00g1nUIakGrPQTywHeAocjHywJvJt0GVlokxSA0qtCySMZm00LxWIn8aCBBANHwxTOXD1XwfW
dJUEqKa7NztlJ/uM75a2BsZf/x6trRvoH36wXSqPliTs3+4w8z59aNCLSkdoot5AVnwLurtIeq3a
sbhCnG43aAMGsayxtGq1l4audjyDGsH3yCZd5hvR0hbjpCAtsMTsExNxadZypQM1OIRrBEuxhNSe
k5a1Spe2tWfiJYwQMzjVLj1sCBYkkmRnh+gREmrmhT5nud4ifcbYpOeltbJqzyLgVz4jWca5sYhi
j4da9QxCpYeV+IOtFCTh/zO6UzHzcyFYPAjP9/ge7TDlSyF1MsZwQ6p2VTVz5hG92giSvU8noFlm
fWqILv/hl9FrK8sE8XMxDJw1wyzpvwtDtmWfqR8uTjyGy+5L1VbRuZ0nS81/4X9i8KTZDJkkiax+
K0gP3+C9vssTjA/8oXZVZnEL2Sh7RZ5G60wALWax3/owdg3De0kSu1MscI5dGy7YqrzLePUIMmHu
EgkCJNcz1a/QNFW1uTBvO1XBEkNi1WCj6UeZCa8NupOzKCpFcsBj6syaDap9kcVB+8UikEofPhBU
OrxjM9z7MDZhHQaIkORXc4wiX8DrI+0FxKRA3s/NcYeWffgUmILJIe1FjrefXHS8A5ICUk/d9vqu
DOm7d2tDIHPzsuQJmniBGQriDR+/WxpWGQFO4RX0e1SRT5sceSSn1nJJCWxpFz7xh+SNCM9qWslW
toG4W70DVsgKp0imGNkAULWb5aGqQNAtByPL0E4x/nA9KsmECVDa1fPHSYaw239T/NutPwR7ipRT
fpYVe4dQ8a9mZFsS/UamIAjKptaKz/gGt1v1NfM7Fe4Ti/w4tAbri0ZJSua9lk+1ooIrKqkBR8FB
bu7DU5dDNgjX2YnyvecCFmTpkvQ2tiwjFdDkIVlaT7ZfmlITAbMSK8sTaPWobOU0sB4i6io6ISuq
mkDdXmJK1cc7m41HeEhx6aOrEpCA1qAPtJckTyftrRKCoC05VcqLg/WOlIWgaDgo8oCcuwpXyz35
Oqa5RiY8xghGZi2fbBHqwpJ4HtQJjy5hknhB1zqSUxOop8nu7XfzHEpYr/bQUjE7i55tPY5uG8pQ
8YvJkv+DNLwPxh8hhsKWfd098fJ9XGUqxSICa0OyK9E7gI3oJcj51T7Wt4yA3YBTpj8DH+bxvc+w
ASSa7xaVAXw86j2rUWNwvihGNfmXFEdU/a3hQCcUXtddMRgSAJ6mYHKwByhX+M7OI59fuL4qsRze
GTHr4m7I89RDhpTbZpf/eDM2+JcJvBG9/+/Yeo8cXACdey5peKD5a0eCdcQmQkpE63vKpap1bi7N
Cu/YSsYOBJk8sNK8sfyKw1VdBBuCtzRCaNLumLkK5puQ4L6Ya3HiXNdBsOfsA/zyXWJw/mzbxx0+
vb2KtQ5mj/f6CauAHWlyy3MaK7YZRgr4fPiOhDn3R43fw3e2kpX9s9888QYUMwKHtYHBeHFQFnaH
D4d+N0ESVCuV1yU5ZHK4cA0/yrmJReYCtjN95qPN4UoiX7s4KWKhAjGPLmVIVZN2y7LEcYi9QIlw
vuHPDzYeHHKM9cUXEHUqyoNTC7bJW552n3Q8KnXyyi9vTwf1UTkLr2TLxdTnD9NyVPNWDFT+Od+5
13hQv/TDLLhszcFfRh/8IqB8qdSD4KL6Vt+U4tQ5KyVGuu2Yi5791v3mNq6vyKWCY3+6xXId6FFT
vOYpPwFGcGJGON779rxzfRrj2IjHsT97buj4rzH6dGB53Yb92MLTL5Ci7NKAz4vC+nBY7Pdfr6p5
9fjY7Zd8Z+wJiBeqQbmvwp9QOT458VEzdfzL12e1GHMX/3q2nCbO15DI8do0GvI6XoUTPJJ20lBb
Yhba83Oh+og2YVhLVYicMInrFMFCW5iXjgafHkbmc+vK07/WlLppswsAfXnGysiF83Kgec8501EY
Wg5C7A3ZvsYrAn8kGeHzw/Q/xXDilX1K2rKKZvOTYGSphH+xBunZjb2aYAyCu2P0yeVpqH1XAIbx
pfA8W/fynyxnOTCEONT79aYmzfTnjFfxLCCg3XPvXI6OpO+5bpb8zF5efZO0ScPLcdVK6kJpjiAT
eVtF5hKpntCosGWqFkRqeWpUe61G72iA7rmMXXID53flqWWZryxZLe07LKBkytJPImFtotcPwaLD
skYChNFfqX5+oUpARaObyYqx/xwsit1S3wqK28Q0cmmlpBhoItx1zzyLLHw8V1lgWGEEtArDyfEn
QcClk93URzu6n5enlu2BKduYNyDu7F6/fbNTIWSynmaJa5s+/GolPYZlNrnK6LMIzNBICHRqKlh6
pcVRT7ZcTfJ/8KxQPvB2n7I3eOgrcgoyzy+7e52Q4EP9xPXXWA1ypimAMH8mDtTArofi1ENLY+T9
gRJERMfniohUhg0B9qm8XCRxRHITh+oY94j2xHLE2ZJFYC75UYI7EhEATx2OeiG3+nERZPJBV+KQ
9JnYv/LieX7HpAxVB98MmGDuT66FJKCh2FsXzg+pNO4NtmnixiFSoxNZZFezve3X+3BXAxd73EHZ
zwcHOu1FTTEjYU4CRFbAdTlU4XMs9Xq+IkSu1o9kKlBTV0C1xAmPpanonmw3j9ybzrlF5kWwDy25
LMsF3gVhS3OcLgvBtjREBHAlt2AslySSmVh8No3IYbncoQN15GW0cHumHSZbirHd2iILKeeF/yVh
86zN8sEt0gBU5t1rLflToclG1ICgroi3iKk37Q9FlApSQ7O3IbAt9R6sVqp5EzgBxe4BItH1arf/
eiRmdKia8zetjrVHK7nWDBuFi3S7HCQXWwcJ9fKDr2QTRF0MaWoQHc32x3QyLcM6PVQAslnDBgTe
YK0a8SdtAgL57itg3TfXbxwe2mscdpcEjVuRZsYZLI9pUdLT0aRkVG6zNUXW+eDgKCVylLyA/uA3
VNitz8326bcoZAxo0IhbB1mkR63DkXmWhnbmODZNE+91D7HT034TuaGU5Knn1kmOhiP0NklFpK2B
X4h0RLAYNMUHZ+RJEewOpEt/mSCORs22mHAr62rxcfwG1l0uLSbMh2V/v+p796V4ibV/7LYlddBE
jQ1g601pXl2+seGGONUBqMwiORo7QFrMO+dV05GuDKcIPxZDm1I8x/nnqH1Thwcwgie0PWd5OL/r
qcutluht7aYUIwYAkEBHb8xeimK3Y8ngBAx4nWwcufYi6F1AEKDZq49sEoyHUZYdg2KYFP6gJhJN
4wq++JlAd6aKRz4BtzeNqTSLYayI7mJmilnNZnqXve1ycjNCndVH7hVOn8XMV+PPje/uKljHe8mA
rWYTsBIo5nOlJmF3brvs1CXQNYo0SkWbDSUBekORP70/xwNWcy73mXA7aXxagoj6oS20aqQHDoyH
nHxXfSoA5HrrovEwARR3Kyal+HpvHhNb85NoPOS2kj3COD7P/bfcVNins4OQPLMF4k5JtH9ZIGOj
dUb87aoRq3v63TinYxCeQVDhYI1DlJ9mvCOZwGkNXg1pwk4xMRzCJhGQieksAB3Q4V+FTw+dz7ib
u1KUnnlbuPShn9kcCo2cdUZgkyJlqvFRBgtt9z2U+44dIlPdw8KBn8HgCA4OyWMunT4e+LU5O5gP
pQA4jWeSOPkEYR37IPeuhkUYS/QFyzUAh1qp5AngfbdMwQ8GM8N/pnSTrWdmSWKlKTNqXw/Znthe
73SlusOfj3TZOxptrBdKK9EjkiC0c4JXUWvmntJBc7w1MB1jZBs/nNKXG2pu8Ei0GWoH88MemqnG
4SLfzqlTkV3eBNCt8Lu8745/QMhD6cJLvtR6ZkWrgRTlpOz7Mb5HbFFrtjtH6ZAlLUWr7EsF7AFV
93yvcDx3j3qtAzCMFX+M2eFQk2HcIa1d7Qwm3JOkztOUrpcBCj/st7k0d3VPfIL3FkW21ukUx1tt
P+SzcT0Ek7n1LMKTkO9dBzwklnolbuSDxG3o6YCLaWZatZsln8ctB0VV7+LdBk/XgwS5XeRuqnWP
7Ia5rTaaRXzvg0yr344LpRIxE+mMOxYdR2sx5fxiWJUIc/Cgh49vNOgOrCnYX3Ac3O4YUXHSCQ5h
LXFuCkmM2piiNigbCd7B9ob3jxYqLFX2t8XunykA7LMlx5XDBD1FmtbyXOzq3eDYRDRBK0Un8e2h
2LBl5giPiOnqlX9NMIfzbhcQhJMtUERTAM4WCeYkq1cVYZQ+sz9JiRgh3ccppQ/deoQwx5LLb4N6
isgpiKv3d+VTrJsmRrLIfEELetY67Lhk+rgFGKrBeTz5IOvQgVQ1hFHqtD3DknI27lckowE/kuHC
z0W/RSfX42qJ7/d4G5hwSCHN31HdJgWN5o3ohy+Mrqq63Sp7fuz3lh+fxelg47T6uaui5WiDtNNS
7GZ1uaJnVh1Z2WCr8lVTL9Pz5mt5RFdtadWIgjHYXOb2ltC15bYYB0U+HTu0XVhyVk0JH/Swqixz
seHyVpYXsGNVgeH8hEzP0iAj6DHiZ/ikdmEO36IGJIkp0IQSHj83sz946lk/PTxK+mIL8yn2xTFQ
yYUq95ipHtiOP6esCm2/9+LLpoavxLm91BCms544w/TIOmBwoqOpXFsqY5GS12S/IQPiJdNvdt/d
lQwMH8BVoJwnUTZQjwbNRE6UPBSVM4jzETLa+5CmASyybwuuIMMabRGmZR5WV/njiHagWVpCk8Eo
cIN+8hQyLeBKlz4lVfcsE/Tc/bgIqP+Uf78Uwm8A0tgetfV4PGR3EAQitENZcALfC6zZ/TTdqHGP
RdN4OqinOmFEC/TlcsAOCyc2ttcgMYzHIrcHP0ppYhwshDNh3PCL9SPTUBjZ0Esy65Sanny7GU2T
CyA2ogGTzIewMlHsfyP8k+6c8QlStNaRlXQ4VBB14s1FdCT6WfckU/Z6jJq39+z8xP0jUaO+vmiR
lWEb7PRtRZvf8Eu2nzc8qMyJtvXSsLNQfBFnabRtAzicvT3ztmw/pEFZHteH+i3tNpbzP7OyyLze
3zJLHjs1fWdvs1vt4uP4TQ83smvE8KVpLGRCU6lSEs7hUcBUYBgkoi1bVMz48T64/1XOz0FYgGQR
/Y80f/NRNMvZTRAqH1ueP1lNya3vohhBk8WvWS4NwofwlyTkvigea2FUuxAiKS8qeHbx2iuRhiqB
QeqEpHghNdO0dWrBdiEwdmeElJn6xdnG0cxq+geTpxdz4HSy/Tk5ivCSN32SWPagnQh+xe+yQdwe
3aJAk5ZQJ5K8YfMZ4HG4eDJ/LDpOo+nqusKEU3G+nEEROHidfIzIjc/RBucPfsP/hQP8i+ddCM+6
aQLZNreciOqWmgf7/VG6rZxx+BB3OixfuhqV/PWiG0xK8pJBpcGlpH67Wv+5t4WYtDWzDbzutA2O
1OT8Txyi+Y2XaV9IgX4G9qFUcS+3c7mTOG42BjjSNsgQJhIb7O0m/KyU6uZuTk7fbKUOWZEk/OJi
oss8eGM2Fot4nFwTby+mIWRjyTuCgrb+G/1Day1Uq2tSgUR9AdbP4sa2ieYbqExRRkRQpB8Wi32F
f1i+MWC821edsYgsYhTH21fvear++MGDCaVYYnkv7XQts8WFnpkjdK7To7Avy3IK8TLnw/yTEj4M
3bOyTs58ufCdqydtUWGt7doCSI7FwoQtZqWsBQS4szkWEWMtMb50VuLOwD5eFZCFwfkbLoCtSLqT
WjnkTreMaSWcOXhnPLPTDIxPSDOF+XLk/HdDNWd80+scCSKYM82bdL3+TGAJcUbCXYlUjFQH2ivl
CeP081mhGI7gfn9CzdOK9OLsh9583Y7kzqm2pPL+kCosQ8pS4kvOcV1Dg/0EvGdaW3YyBNGGV9Ba
Kn6lz+i5uV76W7SG6cyIvfak3Hk/cPRFQq7/t3R4VPPasiEV5N8fUV8z8xCTTUOvP1m4mIr5n6Q8
hH0dO+0+QPcjJqcbj0lfyzLtxAB6R8ZNtqsvj6EC7lLNhDxWG4dne+vsityVGrMgdPVmjdbBvoU8
xpQG+0+nrPA+AZ9coSMWXhxpNzDKi/drDxOrorp53MOnr8in6v/+umZTQ8WyjfPUGzVLJOQjlrvI
mWyfQsvOQOAdKdUJG1lL3ZRXhBczQpA4vDFZ1KbbiTLuSUhSDxhVA0/tMYo5Phd632r/E17df3iK
neKHzsLifMZSPNcCHU04Sn/Tz5GoGEOZsF1TKM0qk4BY3MdoO55IZM80xTTv7Wbbr4EOxztQ324l
ioNwmuKMR2A0iv33ocLbzsaV0mNqIojOBrouBCtlnzfMhX1KanLCgIs9Es6YHYQnzWOa57VGFYoR
lZw7ye6LIu/Pml9ptUIG6x1rq4BWjVhENhpWmbOj/d50A4/wZHBd670ZpYJzehNV97NBZvGlY0qq
ypdBenYCZ4kmRnc35dBwaoprArq3Rnl7kuoMLDnAF0Ale6UFyW5dDiCCyNqGaIq0dVIKGZk1NPJZ
gI1wHuGQn8rOWoO4DjaKSXB0EUndtjB42V3LbYFcfQowP4adeybWPwldlJJhX9Di3yqKUZkRHSYi
0TrjfZ3szsQVkF7cjrE3cursITZmIPNK21KJw7uDYcQdS3eXViQlRzkqYJl4wjYhyXwZAhbe8Xmj
5cx+wktnWOnl0ruOeB8jfO8vMdXBRGxRa4lLC4q0R5CNS0qFjMI3VnEEb9mwMIsxZQtaIw+LrXGW
sRaV7nEyV125YB4+984xMyPOjXE4VSr/UQze7Ob5U3HHdOmzsWrIQZjLLI7iaELx4kyGCFDv26yU
3Gqrii8T/4iuWXi0c5euWJcGWl2nRkC7MpvXtf+fwnXdcgzX8SRuai5+yvwc7ReoiOD6p9WOWdaN
Wb063mTha0niLNJhRVKpqw+t2kCgNCxpxQZMhVrpEhuPhM+XiPeYWW8Gq3Ln5S0wWBYWlDs/9H8L
v8L2wuoYsYQHzML0JPhepk+cuJqZtV5Jx3el4Gw6QidfXGRsTiCr8dBbDpaP8Jzz1xy28sxkG1EZ
frIQ/3EM80hWqSXabDlgOhMRKXihdKcjwcbuI1cD1MoudIDw/G3a33+k3/Ttr3BSZzfnG5KVpIuh
csv5y9En2aZGysNVPvKPK9EvAcAAF/S0K+WMuV8tkb4Q2iER8wnlx6p2rPY3k3RR1XDOTrikiWt3
B8rI7BBxrHVvts8TTOqcp8y1g8TGGhYzlv/sJAlI+ERUGR5yRwPDQXrujOydPYBUJLQZjtAEZ+Hx
Lm/R9jOHUsfoXIopbSbM1SuwEqCsSC5dOIiRXZABohNObcsZQpV0232vz7UjjgrznP5qjtCCDZbw
AcCRHC5nUWhAGkqpSa66PuRMNqHq8pbAzrWzKZa4u3yUB1VQPJ3ip6B792Oeo8KUHz0hLHZH4jfJ
q5WEONYqQuuNVoTed3/fO/g1H2b54FLmme2ExKoVGgPnZHro5py6HosFnaU1oO/+Xul6aDhaa8nR
Bd5SYf+8nMVJnTnkmIuY7ffcZo5HfGLWD5YukJTZx4PwfaiTkgZORprYrbvcOQJCLGJuHFOTXQRT
5huQBjNlUMaTjbj9oOylY2UB51kCJWJsH7Ilgm9dKLyBsnYcBx/1nCni+fiRdSw4c0VQ4A+ZybTs
/8EWLyMdN/skzKgQl2gyKd0Zposhfq1Z/0c4aU3JyMcA1dW6MjCwby6OdSLzp3D37OY7B7bJBXty
bPZziUS+B8ev0DAPWpigF11/uiStUDJH/A0WPhTn39PekfvNyOxjcGojgZZPSax66k6VEedkstLK
E3RYuha/WpM0Q3FQGiieUaBAE9RUC3cGyfI/j8b9ELKzCSGgOwQqQrXna82sVfYgYPeS6X6Vhp/S
P/LLGrdd3Tfu8ZEURjiakMJSlrXABVDsBAyoBweiw1Y0dSswNuyTJfJXPAPUQXGn7lbpBxtkgse1
5vfLeW4vFSR9Jg4j6OyvmzDet4bsXzyPLC1dEM2V6SLeR2mcxaPloHNjTs9Ti4ufucvk6+/408iT
caaTawJjsAzC3r/5n6u34aVNKuK0jRjeIiNBfWPR5lPC1D/rVnucRT3qWJ6nR7EmDyLbTiAa7Us3
736QWP686zrgSVUktjjwiNMOG73vJg/hB143qwWWrmobwEJDJJ97uKtN+vj5PH/usgnTlwAoqrw6
07Xvv0kuKqm/Z7EnV6IkM+krZ9uCHp4SGOb7zm3XLwR3si0Jjj1ePGLS2ibLhP94fmwV8wpUx4Oe
NsX1t1hkhhKrMNfuMmatuKgGTB0/sGuH1GCX22IE5QmCfx3Rlohc2Y1wb3ZEcf236PAHGlq/dnoN
9kNb6B8SJyWDvTmd9VRpiVQeGMib2eUz1U5Ox9KW9JK+22bJZGxvzLhZzG/lOtR9NGiWHAtzSHYs
EUl5cyqWHsk7ZNf/+HlaL+a0sD9/yydxBYM/28CdHAixsrJ9OJk+uEc0QQuCll2bHC7K8CvMNI0h
j6Bu+NjV3YO+rvkiELnKmJ87lLUW47FhI/bJcAwOih26JMDJtgdyuPkmovsYJ1+NILH9ePLSyxPP
xtZjyL0ckpaDrAONeyH2RZ7jAVr4SYqqY2acMcpgKz8RNx+CDIayqCOL7fy1OUuZmiQAkq+MVlKO
vNX2CV/5ZCt6uTxn2kmD/Z2hVDIuqZNTeB5W00/T/l3bOcZarlWyJTm2TXMMgtvrgqsGF+JgnkGX
Pqc5eGFs1oN/gErzQQOy+9BOOtmQX9SN3qL/eY/ohOQOhR8yQVRLaxBF4hgq8n8lYha+C9FfGQzp
5PFsyVVklPhSnzixctVpG7eZUh2AimCb6/CkutuP/3AzZYhDg/XOwK9IhnXO30vfwJWlmnKd2dNy
fHN9FWGbCzp1GvANeYYRIQlb961JOUJbMoEV/IL6sKAU6H6zq7Nb9s4ueIHKDcTHo5UYi/grrgQg
q8pqAf++etejTCz/Hn6nfL2e4B3v46hjYn1p5L0o3pbHBG+AcejW6IXnAGFICUlDgcqJ1pR97Yuu
pKjUNaB3ip6aCtg1CRP0hxPFfie9NvvUCcJJ0CZ3TZvxooab5Or9/g4HxVBLdeIHOqp+fsPcu7oI
PfjP3KFvLuOa6ak8R/bA9a0KXxiyoPvV9a2EyxTMwoEyBnXelAmd2ir2EUquW3EnvOtU7PF6s0aW
nIo8nCmcWAwhAfUNOLKEaaDycglMrjmWV2WL9Vu8ClRSwFhLc5jHMc7aUxtn3ya++LLsAogEnXvQ
1+DnXznHBtZvzycTeGAKxURSYueb8sstrbPHJxADNHu1F0ToC7seHze71+ft0AloWqFORBsLDOlu
G0a/6B0Z5Vbonmhq0Ci0dYp5ma+bpBGG+93Xrh42k2d7oy1MGoB+UEs1UjZgir8dEKy9C/EgFQg8
I/GSX+r/lzYoJv+F5h4K6qS9ii37PZTC782gIJPhKdldoGEMVh8gsN9H8/1sqxmRyW2fZSgKmhhe
2VlVD/Cv9K4Kq2YLh4mcO0Gld4djAiq0VJW6WX2B474bRC88lzUK4ZDy1Xs0BCUKwiRQ2bmQG6nV
mQ9a5t/b8Cj5Cn0Zczm4IEj8TWUBuprFF8C8meyeDJ8tpS66novU0cWMFJlut0QougFlN9DtNTFk
Fv0P1yMpkvlH9vQWnvMANR2/XV8ydzlDTt3oMMMMAbhy/4pdcMzamSU4TEHigeyWgQB+r16FHQfp
inuigR6qiFarK8gsbeeWBwPw3qSN9H2j9KIm4vTpz9xAai6wzRU4Con2Ws+N8aLWlPUkSDZGeDTv
0XC+0K5d2beUnTH/LRxhTMMF6eg82vxRBy2zjBep6Ilu99HaQhUTGoQMP1Qene2VuWtYgfYg0P4z
EVPfwXnwivY8gFB5K4g0d6Bq9+MSkM8FSLaCumicrxNSxJbs/JBeS3F8A8uYpPPf6isTMTjlwgT2
TWmDdbAfuguERV8v5d+Mza1TzTKkjQkwMG48O3Kbb6ZeGFqat49U8qnQVNAsJeiMcXq44XCMf5MZ
wEUYo4dPZ22Q2yx0/sRdWOk9urg5H68AxlpbTT2LFdV7s8Q3/bzx1BZ8heONQg/aU3gZzUpZ4is/
a8aopgljlujfzDD6ST46ZzNklIwPb46r2pEjYuAs3veXO723IGk/RVAFK7WwySr2O6AXDhBSP09U
YQN4Op6Bv4mQ09FhbnhsL1Q9fnAYfzfaYbj1HNY0uM8t+82FY/auY+o80WyDoeMwxLGvejPSRD1q
FPe+QuMawhOr7NGSmiyt2oyPp9a9s7NujFGAiyTU1Y71J5hVrS8ONXRToQ4AVN/3ka3x0m+QQI05
w9WLCG8nP3elDU/NjEVwpQh5mdS/lmHAsDdwtdnithUIHzhdE6ZaGwq8JaUmWJhNaaGv3E6KxTl3
DgQ4v4hZGEw3KCcUtPbbzsrUyEwpEBIyIamu+phx+MiKb9SpQI7TE7DFfaXzkhFn6GC7tZAmBx/3
tiJqfLudLIcqOu99uXU5O54RRTpGXS5Nqsri7KDJeB7xnHeOoDJjiJ9MzJWrjQN6RBEuAYgzEj36
oPZJH49HZcHML6pQYD5rlfm2hW5I1VjF+k32EdsiNKa2ideckn5TqSK5B2A65iD3amlg5h5MQtgr
ufUzr0YC4qDOwn5jmIYq54g/7/6juSSXOlg486/y4es+KCasaHi4l4EDyshNHEfUmqNRXHhOvKM1
xoxtxNhDzy6gUqnue6iGdb2H2H5rFacs7ZkFwtf78lVG/6NymNKJwaENlrMmRXaV6Wc0Joqkk+kF
O0Kbo1gvkhh7A4MU4C7/nT6mIpUGHvTEaC2dZAYfOEIVy4iYBr0VPZMNtOGOENx5eAOIs08OHez2
i5MF3gUHg90agEOXIHXe8YvKqW024nDY3OWS5RThCDAjl96m7KhC1586795zx2R1Zo8nFlr/9XYk
mHdyIicKRFPoFk+U57QYZQFgb+kuXU/exWQwvitBRES+1aPROwuZufLrZFEALtZt5AH6nRTxgjeJ
p5ef4vhyJLdYsounacSQg4NSKeEoHCU3QoUvP3SaWMslVSG+MMPtW6TFrOl05V10H0kUo9Llpulz
RS6bCSezfuk6dWFINfeMZtF9mWpXk2NCld1SQJX3W4Zdr3rT+cNzEqm5SDdES7d3rVCicXms8x32
0dyJi6LjFxofheFRSBnvYtnI9ytQDE6gEAE/UnPIANc1nGz3zF0oSwguMiaoBlg8Mj2OxbH6kzwO
Q3yRRzz9QhEqsQccNwx2SKJrLrILmlevb0sxRbsAMOfMm5r3io6NDnyNv2o8+B8dH11v6pq4je5x
Tl9Nx/BzYc+2txQDbSiUVhSxcpabjRyc3WIoNejpoCVznojHKJkVy5Pq1mfhfcZpefl0F9IIiUUd
YLnwevD1Dzl3LudQI9RiE8epyGDzVsw7SxdZbrzO++h5FWb2Izlmo2VaftkdItI10s9tZtmC2HZ5
+m3D8XQC1hkcybc1G/kme9oigs1RnM8dNIXUTxCu8VqsXr44jduTX97Eir32Zn/h35sWQWtJPU7n
N0oNhTUORkuBMa/vP20cpi18DJyW2M7FZKxpGlNjxOprShNgHXxZBp07wWqVyWxwFJhJ8HPeMxg4
d50mHwcfBS2gjIhaOY3dWTt9d2mpIGCijiVeHrWNS7WXAIWt3g+XJzxFD0snXuMzldbRcQ29hn2l
5/M/7PBCGUA4bcOJzQqz66q92fO/UsTLWdU68iuO1Wpoz4gMQIb4ff9BTlSnSAtN9/TXILKVTo2b
wE7DoPg/6iyeXz9nUB+TB6wNOfP+cKGCke4r5vOndxjrvXkwCgR0BntVTwUzFOWyQnJ/9awndmh1
WrG+liQxGRD884EAwUAQErcwwGa7rGatWDEL7/3omGPg8xLkmTss7I7Gw6QKLX9+jqEdqLIJ6MOQ
XOOXlNsZDEtbCKj4jSmuPF3YONPze9gfjTDbgv5C7mNeiut8VyDlVeDmGX3L8X5CY1nEgGcShaM+
MvRu4mxzBEUABL40mjtle4sSqm8JaCP6buaCHmaNqF4xOpPKkGs3idCUVqG0zP3Py2wzX8m262jK
QAc3CKpWZSV4oy9NHQokQO/wgXl/BK2DGABwGp0FgwEXpRJ6ZSu2DCp1qUXXtqnBcE9TjOLQbJcG
A6RdMxkeWb/gOoUau0676SVFQ8OsIDG8u4PFwt5a113pHNBPFALGLdOipOM9eK4K5esFX4sHG8mI
x6yT8cf4VIXOV17jebclc38p+l7tRg9/iUnX9Lw3n49LYincdgysAzjfCZ90KSQublPWgkzfsaqV
DxNtLgr1CdeV4h8LtbO0BGQIT4J37WF/t8Ji72YlafVTmvAUsTQrZrEAMdX3Jda7Zh5G+ulSWj3y
mI6moU7WVOaNNBpL1FC/picWObhSTF/A7kJc+MrYVEuZKBnncHnS1DRrLz/Tq+00Mo66UoG76Byk
YH8rI778bv9MAhqE1YzI9fZFBmgTHChVtSDYFNs/KWy5aHdKC1n0Z3cBNfWDt0jam0fYKLvgsK21
Cs8iKPKewKv5j6wQ3x9rXPh45JO5cF491bv7ob2Ini0bXb8o/Bg33hle+zlSqTX1CoenvY/iemPv
a4o6XNJsQGxnE73/47Jdqnutq7keVCCBaRn2un8cGjDRrSIHMwSUvWvyVl2QZGvH4YCT60LfTlmR
YX6Za0djO+Dy1RtbndIkvuZPvSF4D12Ac/PGhHQmEqeG2gzacjJi0Rnr4gKK6Cb8HDTPjinF5fDw
x1yi5HgrYJABIBlmPB7UiQ1vP6Hqcbgr4A24are0HGlSKCWOASkFG5EdRyp3s4d9HhwPpQ4duFdL
ec8e1ZPIRBceXeluQm7N/IaOnN/EHSqoKlseorVRbEKZ7QVjjcN4su5lCI/GGrfH1sP37cRaZu9Y
x0A6UqH27fyW81ujN7LiNb6myB5K6ksF7tUIFYaobk2UMje/SrEeIqhPiFi1FaTNs4fwYBqDJNJx
zr3K41h9M9aH2c1jdzsVDCG2qfX9j0UwjElD2dYF3Z5H95GwKPpRZSwazPAc/mufEuP/CtYAMJNh
Ut3/3zyewXfur6Mmg+fDMlWuABIBh0DKv3Aac1kB0gawsO9xpC8QNgsUb20md/0/nbc82v3pPpst
z/94YWOsbvfztjaaN3BbHNEwG5J0kk5XSyN6xzWa1dBt+xStn5sR+alOu0QVLlw71G0oDTB6LO2/
f521KWzMxfH9vnDPnlyvOfhB3e73AgtdSKOc6fEb/yxLj0o7RS3aXfyjv05+jRb8lcRswt2quE3j
ty7xgE0E15mwyvX10Vkmiaqpsa3fKVX90DI8FPkLgm6BK/nPlSFsz42n9w4/0b2zDJUjxl4pPnrA
6JBFpan4H0GW7PYp8Cw4+mkcCQ4hF10Lg5ZTIBZYMtUtR9Uc124gVPsIrBIYgdVkbhlh1mR+xZxM
BMD1W0xDUeEvks7TUwH4hW7rKSKHec80wJsN5kb4mOCxo6hYtfmWSykEysx28pmk8vXbVeZhWBLj
i/dPmRbMGTN4aE3kiMJib//pnF0oY1ARexEodUoY0i3RJGhjMM+NDnoAt+8J4lUIH4iEg9Bq6L6b
5Kc1RunDolSAl0bomoxHLiTPmYrhMtkFNchUPWkLQa+RuLNfszZKttbieFf91GzC3cOE1JgW3/1i
f7hbzAmrRSCwI8RsEddJyinQuUgJR6I43mcmkLo1T5hTlXWYrGcxIKXdwzfvmas8Ao0JYpA1t6Kk
+kwkIpqI7OC3Fa6DmiMsgfOFrvMiaMCye0T6id0V5vmy/TnBMvBh4ChPbuvUrYFbZVotVceHdoCP
+qpEgbuTJ7ZrIL8a20MbjFnUiErzkZTEpzSCVn18NCHWoTEFbKvfI8OFO/kWFLqKQfZp+rSOeW7/
ukqJtg1MwrRjPdYz63NVil1ru4v+dvVk5uiQPrW3htStJY96vlM5Ll3/2qj8bn871CrCrDSTOU4m
e0js6QBYQKtdGq/2H2cPREtKr9BDVniXTkzgkVOrS/ympQj4hQLhqtNxN0Sh2lCs88yl46g68/V9
8FNcwzt52ykQum/L6bFgrUyDwzZfPfPnGK7w8aKJsAzJ3vWUt0f9fqgfmL3AzXdz0QiT2bdJKvfg
uejov2SxB698juPc/6wJJSkilcwqX1WkSamnhbWQNpyxtxJGLToizxjsud1l28EGRUrIZ67cRuJl
Qy+qI/Wp6LbMMg1T7TG1Ssz7R818rQexUD8pmGklD5n7n8vO5+ZWq7u0q215Ho9jQn4VhUxFZg37
x8Sz+lllhScpIVJhAHREJ19/RI6ZLHA8Wf7py1KZOZjhS+b0iIwOBsMrIhjr8g5GoTqt4Te7epfl
suNBKNssANQtytA8oCafyUx3wQOi/9hEAV1yi8nKBRQvjw6KMHf6M2xrzBPPiezGDA2sBuJOoq6P
eQ0Tm7XhYC3UR0TNYVnGj71SF95z0T9eUBx7q4xF69UcGh/o8wV7UQIkODRdB0jxZoV3BXV2vtVY
6kd+ulUAOYFJ1sDZ4t3rGLIxAZ+OfXe3oAFFynUM5AN0a0is/deSUePBuH05L+xSOtrAjO2Czdam
AhT8TKCxrT1+Wbbna5McQZ0IbTQrAOcf7m6cT9tjbnHb/ZN456njhmS+u2TGNxZeCCA26vqyl8Hf
SjnnO0dUziywiwMJW/0FoNSDO3knnrmoL4OFvO43lQwAgRWYJKg1+SvQdBgtBNQjdRTgGu+MdWCw
zpLjECYQZSNnoINzeD3NKZEIrgWNlg9ujL7g4n907LACfeS8xqllqxeyky7VlXAUqt5iwfFk2K5d
7+st7YyXWZ4RUyjUnoD1TVt3AILDasNSmBBVEOEPm6u4O5JSWziPeqUqxh6DqRV7huxnybvTKaTN
xJTsi1JwE/Fg8pMsa6ORBMUr/NOnlYBtCok3pMwgJ8uJM5974r6M8M5UjCOx8LHia+io+mdBikE4
Xi34lWi6LBdC5GF5Wj5D5m1t1D5HymOVkfSbacTDj6jYwbky1ZnMEMpF+CIPNEK+fVVBScEkhjw5
YdUu7ZpBkhsbWHehEtBKWSxfzYEAGLmTkbqezlycrAf3Rfd2CtHTqtsGyfmbrG0cq0tN/Rt/l57Q
/rA89bd4Jf56YFgz+OTcyHQHUubTJyowq8BHRVagzMaFOvvBgQMoOhOghJpxI/hkenID9usFuMhT
gxVsG4+Rkkvq1ym7KH9l+uuGCpz34xsoghK45cK1kLKi+UfjW2ndngYtfhmg9wKUTCqdWac37fxg
LN7WIoyoY8+G7HVXZEn0l3RDbxRKUYBOrv7z1EatswgPPHr8h6EBWh9lr7kNW0T4wdNTwBZ9xyI+
Bj/sznxtqILH6djREnyqeaqT8j2DbZdjQKfmTDU6fFoxyjfkQtkCDAJW186fjYqsi/gxYeCMP3dV
3WkyBDHA2oH2CrQcO+VKbqqYnVcBzG5yshzNufE3a+Lq90sKb8QGCL3s3bTZHMybC+H/BeZV4I0U
RHh6F09jXGTTqvRo08G5IrwcwgTDAsBIrIxyIojj8CdhCnMetGHqF6zMEhAqU2zHsRa6zk0XSxx6
DkrUc8cX5nApR2v4vh1hkm0AGFL7i2rorQrim1LpI/lNBp6Htl93mGRRtUKi/R5YaRiKiI9IhSWP
928/SkE00iaIWO7MGEgMKydABaMY/qGQ1bG2gLrc2J3tdsHcG6vL7/G5YpdMzCrkj68nALC7K/CF
2nt/ypCfp99EESJLlBgnaALpi+qM+QMGU0ErDJ2LNAtb7gzU2W2V19gUqVwllb6FgQdA8kuFDmrb
K+y72fpahhSFVAejGeEkgwrOo6imxD3GXp4byNNA1EXGpNX5ClAuCuIDHRGYi9RinHIO+cXPEBNt
JKq0KFxbQEtMi4DDw8FEKVxBmnLhImy7/jhPMCIwscFKJPIfxkjyqcwV3yJnA1bcrhqS/Yi4hIbp
Esmz4Hi5HSVnMRCjFz3f+8EqfRCrbASzEZyHgpxAZ+ND1pvTCMWE6NBzWdMzzI0WH1UyPOONuone
EEkB6Z2TT+DEd6tg5QfizJPby3X6OZA+NHRt8hmHt8nZ9BfX2+PUgxpw5oXP7VeAz4o40CDT8TtX
S3Zn8xJICKaQIYNtmBN8vJX/ouhEQ8kxfGw4i1LW9qqQiUaNsdlubffml8STHfCWBFZGlo142sdW
6YLAp3Ux22tbULmRY1aquAKkQq67XwKljU9M3FLWdgGzlyZgeYclTonUy8QpR25tMRveGP4tVPox
jG4gbHz4LrZJ74WrKL5jfohxcbabq9H6CM0YDCUEhk8TVCRPVm6EXmf6Oxn7db4AmXwfekfVDEC5
Ye/LHnBKzTW9peExmLSnNGqVWCdZQ8GKFbqVV8uvWxQLn+t5z+iYdUC1ruwM39VyXM2/t9LJf2jw
yiD8LrDEwlcfbovXnIuFVK7DQGugqh3Kx8NH6ikjiMeiNNJF6hfmcRVY1rHMIS04SgW+AlggEKQh
p8uCMyQ6kVwOII68RFsTVEgtny9ns+B4nSRwb/Z/PTa/wm5dW+DlxAx5/0XTacykQBOCaTnkfboY
xb5LoPbq0SpowoS8V2Jb7a1BZdu3OlwV6YN78xvZntrjU8F9iKz/QKgjvyLIVJzlDEA+q2L6ZUKS
V59x52xA5p/O9Ghzx8bWSzLaEOUDWB4WU2ulNSia5zNT1GULu1hOrmoCETMbCZzADwSy0fZXq/ga
bbkL1Y3+PEx74rxlyzg4vzB/fdwVPjJompUGllTwZEWw7DQx10nyj9ykSF0/JGrUxDPaisi5gS5/
soMnXzP5MViXeNh6EVAE8tal/0yxUcx5hl4Fry66iPJMmrDKeV4AU/JD2J0tR3qieak4QTvWu+a+
EHbKbRAi5ybs+zr4M258KS06UG+Dy6dmquv/ADDOmu5KD81yrNxotciLFjZH1Z8HHUM4pHvd2aqS
zrQ9cnslwkVwQuqaW+Occa64pMyJ3rSu4LtJ/PRTiwSoBhiWzD9bmVwm/hgNihlBcMGhnLo1YziI
+lg3PNrk3nBz5r6GMDK6kXvuFUdkrfUTGe55+m2wSrw50+nYGT5udjWLuovMfLkXHnKmfbwNL4/A
4SwIpkq/nrU0vsK9Xj43RnOfUd5FBg3rdsS++sebcQfmYu11QX5i3Ci8F3mIAcxyXd0eyz/RwtxK
eHRR9ldWOGNbyrbCpLG2GNH8tx72ZdpgYlWBp/lmx8B2TjJeo+4vbq2FCS/irP4/VfJRPKDijJhv
80NUlTMPioHbrijNASozMZPMfVPDb+wQGnCHwWFW261bRh15v6QHVLhoMWH83FkOAnzjfZOqxgvx
FBT18FEiBUslsyo3xEgiPzeHBBQnyARHSNcC3MH4/+P14UuIJvPkQBJ8fgqBZ/2M8nK2YXsiHziv
5vgTRspqvZBZ1ziX9INq2QAWBREp7inIsw2z0zi4igqdZNyVno9e1DqstX5gwtOrtuodjOh2CyFc
ZT2nywNnS3bDUYI4baXY/6N6pbLOxL7eYAflPvSWypCJh6MDFH3D9o023TNmqE59YXlowILENd+c
qp6YB/C2RVYNK00yuRjvnQhqxphe8HnXtKWSlF0xMYZViWazeoH7Bs59kXEYpkShZTQC0S5E2yjr
jqaRxrulUn/81LVCSvr8pDJZNGe43/omoBPbfp6Mm8MDaQy0K5q2HVozy+uGwweTW5ZSisWEt4sF
PeBpA34GaRYS0uMlbYZTw4h2xYq/cT4CZn6GZeI4uMHDbhzt3ZQuGABUTvUDcnhg7P+qDAdP+EnO
vaVVnwhHoy9VGTl7huCixE+k+nVm92LdgLFaN1jSx2mAlL8sO4ISWBkx1xivT7UN6d+vWsKBA1DD
3fCIcU3VazUOmci6+gGNtVnmqtk0M2JIwNGds0CWh0v8NLlUkZH2r5u5BWjy/GvXq0IdppvzQ8ki
al5iVZ/xVbXXINV/IRoT1L16xQRl3X51Z8+JQcbBOdXWHJY+rhwXnKuGL/ScZJbxDgjq29A3f9G0
ei9v0njL4JKYqWtQE8oNjXZPrtcW14ympYnVNaZhlDhd5yycivR2LqW+3jzoIaXUbPZF+B+hjeLv
Um2gH/dy72RbYBf35M9UnVcZcyvI5shOcN0fmGkBmfS2dTLZq5DJzQpP0LUDFX+i8ZsozikyjcnL
slhdrS6TmaTcE7D2pB90ZSwk6gSWtM7qu6Ir3DJjix3fv6L4rMWnZ8BqF4DlDFlCHLZIIaaQ13Rk
cK++E5dnVQxGcwOotCzjyz3NgdR2Lm8+5ThFAhXw7Ps3g6D9Oi6VG4qwrnUqqzLdvyss3j09UMlU
38bwebDphHjx3IdL6/m+SBt0xMiL8qV1kZE9/0prVH7KYmnMhYiMCVwOM/brAVDw+ppQlBDp43N9
mORYz2MX/0VJej7xbaAWy8x/yKu1Zpf5HfPpV32VJFMJSMHchEMWUTHGigRFhove9/mNbANinmOi
v/Nppgls/OLITjxdAd+f+2hfe/7X3X4ZyRs5osTBehc5J1vpeO+KW15OXARiazBl4qeV62VupY3D
LKDTM5GoBxHylqq69m/OfDolj1LNK90ir5KLo/PiWRwNkjMKM9sHzYKm3xZNEUXT/jxtW9ZG2Zd1
pcLKmVb1Gm5At6KfVw2W7f675OdVAGBcfABKbOj2bw+Mgs3FKachfLZjuBlsij1icZvT9qwtkt9K
Ra9dLs6gJaCV2l5wdvLfXOHO1cZL6SAhdoZoeJ0pYiZh64nCiJoUi8P6ykcyTNXHRGWhl+Y16/il
F1CieQdvGj+u2I/j049BKN54Pi0dqJ27joH5KfRyFMOE2Fy/n5mK3s8KTfB2AAavPAj4ljwJXl2O
4ycYZBAKvsV0uEBaqvm3ZsKBRi2lub0OF1FA5AXMfqsx64f+klhX725BMFieBqL6alippmSQaJZN
RhU2WVoOecLuaZTNTBuPJgTPA4FaQ86unthWAgb5V4UEvpRHeqRdz0s3QQCY7CAWK2IaryGEEq5u
7VDaCqxD2rgX8k+A7POxpyFGitAkCMfs1aeP66FCDl244+19FZHEsRToPVr08aRqm0yM+nmwOQKF
wxp1uLZrfrqyctjVm4nhy4A7pV1+4s/ZcolA/yz9+g0bg+BZhjqTgf6eQAW0TqfcyLXLCmbWeIhn
wUS+kxQVvGRxhykoN3R78zChhncvyKAm5NPQtLxNqradrtKq4oH3zntio58XTMULWtVFNpVQt6St
BP4utHt+QM2kVS0enUA2siNDF4FmatkqzE4T0OgxXSONPw91FZ7Wq5b7D0g7f1RNRqerU9kYe7gi
iQ87ecV0fZKbW48RVzqUriCLJ2omcbo5C+K9heXdAJ7KeExru2JfFJggCMmTBY6w/pkgU6wfrz+6
NVTdIwSFifvkLjH33enI+5z3ecoS2iARH3H7XojqTGswaeFAdIcCjVtlpdery8mkNMH7Mnw0bNOW
0T1Q7QckJ8Acg6hF1RwgSOznnwl4F7iPvr62DhPPqo+8qYpdAT+IlbGNLJcnmXgywUZ4JyambT7n
6Rl1XtuEElAxUjEKIfQlV1yLzRNIU5O0g0jOcE/hQUKNmZcCyyyG0fZcv38Bhb23VJW58dzr7Nzg
zAQbTD79lRhFuhk8B0B1dImTAtg0oXJWB6tBrr6QIOI12GMmc0LKPHc2XSkK9ZciHCX9/FgodJu+
fkNtQiMRgonzHDTtwZvxbVV4UhmVnNhC9YvISQ4Dy6tbDQlvAADN3IHDFe0ZucxPfITDXY0rnBXu
R2dTo/OyfI48zNM+YgtBODGlQHrwsPXRkKQS+5Y/7vAYgudy8Ic5OVQmjXSxwCwIFSNHN+9oA04/
rnR4qSDujOBBEuYJ+x7zWVV3xOIJfkOsCNgqvlhp6gzWw6WbVYK5x2bykp60DdkuRTe2SPAscWZa
QacmnvpUjRASv4dWmGPIHQDDb/vCLYccbNyAHI+ZEGlhoV6E17SdNJbmIMe2m8VT1QFYCPGiPvFg
xX2PvH2hMz4iDdC+g737wQhH+q+rhgImXY3TapvoRtwxTftTKq0js9r8xoC9imLsJcnfZdxzJBaY
5+vbGrnw5ScMUr1lvGeDc0GRQUKYszvPlxyJy6YMvdRKn3FBn2izyOWmNaasje8I9r1LzNj0t/Wc
KUl1+fjKABW+pk9u80weTAR1IsK1ECnBj6twvZV0Y+WyW1Gn7yBYmLflIE+LpEeFSt5CGse9hhWs
YPlfTsiPisW+OUtRxGc7tgbBZTguBW5LC+hvbuGnEM3M7qIVQvon1Xi3Clj1AvVjMC6BECe8Vjsf
HOC4kqla6H4oywtpCNRlls6yw5dR33RaUZtxRBbXAXSD5v79F8uIEr22t2mmNhvkR56iKnlJX1YG
pdatZW2fnH5s1nUX7vMN8A2trre60q3GB1wA7YofR3Fk2WIlEPdGT10xmTZKnbz1QeD8TnkIZ/9H
nNM53WunajAx50giBdNZfYHjr8ljuiFesvPivgcJpB+n84/gtCdTAcTIxc7GDjmKgh2HIMIE3FkK
tjbJGm7JUeALfKxDvD3pdIFgNJmnAFIB1K0yD3Zxvj5Lg2m7P8G6I5FYodw3LshJBSRdvsAZkDOO
9sfeJd7iuD8Fgw6v7BBoNM5CtLXfiaFnz4uFdcmcvY5j4LtdlRalGztQXIEMXi1MZ05kP384fqNp
gsCDPAkZmgntOW4BFth/6dF3tgwa95h3VkQuhVme0yt7fDUxxUvKCKCw+jPm4eTE7hkGx1laTd6F
MDV8pcitCCqTfGn5xzeWzGCxkP1PBoEN9+RTAuf4MPcPgfk6skhrEFhT6W/0OStmkETQsrI3yYMd
87eKHOoHUOwAoHSZaitSaZz895NQfNb61FYYkRY73pa0ktGuvVxhe+vj/BgjyumwDmmsgpGbWeL+
ZimNiZOWzfCkR7WIX3WRi4Oa8R5Ux0kDR5VL5akBfD3504IqSAddxVZ+AhOL1HlBayMq2YPupFc8
3/nL6cbpYrAM/o07w/K2//CCiqyJAVI5U+kRdqw5kyTHOwJ/x+QLvU5+jLtoj3Mtw9POQlZVF4TN
JzKvN3M+J45hK2DSWSzAC+osBuH2Ij/U6KY+2cE0XId7A9OTeS7/KkOuSxx79kBQnJrA0v7BfqvE
8zhEalQ2tL8W9fKaXRX6vtiGC+iWCYQmgh5DW741wP9GG2HFws7MEbuVw7D1dreSBKno91nKAaf8
SGxlLcULvAq4iKG8R4dHW2j2huhYC/ccd45vbncYQ8cKsTzJ8xPPgXqbiXacOzLDjfR5AmVHKOUt
GTgrVSwx72rkEROCui4wfRExFgm3yWmqcA+y4o5lOXwPVW9LQU5P+df37jNWCLaomYUOWW1WSvFc
bsbZ7DShywBKkZq2PmC9OpV1grWj33zj2am+VAKbQI2JeyRqISmLo8YyA9LJijz+lx6oVzRXN7oK
C9DRqhinBXl/Cs2YpyQ7MKEQlA1XflgIdFyKjbwJQ4FN3lUE9578cAf8s2L8EP11KNCz41jXl9e7
ayo2EQh3BXeVV5/N0MZqn4VGR49LPD148uPEjrNNrfy4kUa1EGXQ+o4eyA2Y+hP5b5rcZL5YIf0w
4WOMdxC9tA+G9VJFMS29//xQWq8PIcyTuVH5SW+OEpmOx2sxBefEagzT/6J4nIf8YxrtCpA2i0BZ
4ts7cvwvJUxU8am3/jz7W9HgqGtdnpQ/p6949Y1R2mjtXag3OC+e0rtjVOKTthloE/1E/EawCkOs
321zUy2F3SxSmkJv6lxTFDESjgo/1mDjKcHb+nl5sZY4amfbcHajIxqCKSrNlRHjIG5+XlwpnwQn
cKOLPwpO0azz9qRBm6teTKCXhbfIr2gLtei8PenAz/bnHKV171WXDpKbyVEu1QjOQ3K9CIjmi/cy
QS9x1iphnnSg6rTgz6lDlV4cTp/YRl4i+bfuGiqDoN2DNqauUkvsfCw3jcJxpmFvG9DKFK0taXUn
5rBeLYWcFVAS8VNAix1dWS1lN/b91NURBOwIrb+nVC8Br+1H41O5hiDbeqDGLuZuxWII7md73bQT
6qq2OcLpertVXToObKJqAxMfzV87Nb2rj4vxyVrLLhNMHdmtMlobfHVpBs3CI/90616LJSvp/1KV
ujBX6vHO1bwi0cGj9IE5ajvgBs0ZWz9wFT1lwSIcemCvbeDYF0LHAep5UbsyT7hYroIog1KSfOcT
dDOZ+2SLMgQFf6mapo/i5xpeiq5WsXD7P0hvwgM3kcN2isbuDuMhthwzzQ8Nxg566oKzaTUeNK+C
cwDP80bvyAF87mI6HSYOmyUny/NdyA/Z0kS6uP0NflSh8X4jJQDBmL3R+eA4YkbCKnTlI338GuZX
DQmDpmMfmiCF7g7diG346afWE6zJrsJrWbqydj+uptnlf5RYFlNtTFUMtcJ/ufk9/uQ3SaVqCSbN
8px3eu8vx9roY+YWtQIdJ+kP8QXLYx4mMP3VExYvqT/btXCCaGq/GVjzcPP30URCMon20VjXrZGI
09wwitUroI9O4cJvguD4ZD+jZav6lU/aZGSYczT5fMFJDm1hvyN1EWn4Xo4hxLpkqzU2VRcznn60
vO+9JC2BGeJZG/zcXGXMc0UXStM89KWmNeZgDyCu3h0tv8TcUAUaoLrn2hvMOdpHk4/Rkh9UnBau
ujoCuSFKprIDnmLaF8Dyabhey6goAZrd+z+j8i9K+3wh9RQAwm5VA/awRzMuCk65pqnjy9IDXVPP
AdFr/QRBrHiG0756f23Avfb0nSh9ggbOn9jfu98z4WunE+p4m7CcFSdE6u7xEv6NMv4U2gUp2H3a
1V3elYpck2B4bsKgZVFIxfVMjTdbTdYFzbnXo0NYRWmc1laTqT98awnGYZUcsQ2rmrRK6FxcAeMk
HAF+E2D63mX+uxhTvvlRAF3v1CEtuVTLizZ3NJJ/wDMIe5qoXEC8ROIVcn9vw8l8PL6eBniSbu0u
IJEf5cGcHuc9yfIV0dnDUHjaEweIFE5kxNlY8+KyF0bGSTc+kmqU+uWxTJlENvE55YM+X8tV2ZRX
IcBKNJco9WJPjWjWVxphlq+qR56Cs/RZYpEOjV5AJOZSVhbK7khjdWp6jMx1b/xPaQzfxe0xwn2A
qSIH/r+SpaSE84Nbg0lDQj3KFcoSHOJUMYVVkMfS18f+vlxFbGW2AilPuQpE3Z7DUBp7Fh6l2AdL
nIC46fAHX9ARgtpLE6Sm+tFEqqq0rEcKI1R2+g9VYQ0ipsn7jsHajlmYung1B7WhtDw9JQ6VxUjf
zNE7gj3tRR+OY/APJPFJ1yY8n+JAWIT4Z+m5fhrKbMhFO5x1AD0O0E4dFz7XhFL2swqqmxirKSzS
D5leAsucVypo6+8Sti6WVVtwXEDK8Y48DKV8sp879YwJ8qpdAJxHMFj+aejzcsvzQDbwUIPuCGBH
VZ7caN5uCOp8lV2zKJ1kMu9+W3e231fy0icyC9pVEuDwOFwfjwpPJxM1gCuqLhxwSb9MqmxJAIj4
Dm432tm5nDdMWogI5RA9ceLpGNb0VWgwVbyZXM69OG4kR7LOXoihRtIIlVrF+gxaIbkPSyRJQA2j
F3uDUZ/55pVe47hJJZplX4O29RgWkyDLnAIAPD2zBi70C1SJZcptWOW0K5wuTEw5VN39BLJjdNsg
SMNXJulZtKe1O+F5MB+8Sgy9N1ouNGOpEpWK3Tj4E9Ks8+StGYbduoZo1aZlAAzL8G9MizPF0jV1
62p9JTUozqTfmI4I1U/+E7YD/xrO22IeN/D61dMixdXy7tihqoIXKcHWpYBXrrF0D9aTjFrm/8ip
CkFqeHTXY5DJbJQimfDzz2WnXWPaB9DEi7GuycgcP/pHVMIOrSpr5eF0vVIA5c0n1t+DnnAmUgdU
sdxHwwjE9clwzdoWGy/IkxNT/gT8h2eP4KdvecNgavAjzd4H6bkeu52ZabE5swC/r0q7j8ZaEzsX
hhOMp6cakTsYaQwKhLLzZMY1o9Jo8FKwHrrQMjQs1wR/usrYpYFjWhu4vl4V3u1qsrBc/GVzhmB6
zmPYZdhXT5kdJdD5NGNUcuGbnJWiGyONE/Tyn0Rd7VgHUMZXjkOHdob8GUXbGuHxW63rSruEGbNZ
PxL+r2gHoD7ifvdCBYjX/mk+Sedx0bsb+W1/slVnjpYLuu/pKQtOjbHWvL/+i+P+yCPrSNCtf7sE
DKKPREWUoY9xfZwON2G1krbYiRMxqoajTIS+nSLdvDRu2CjHMkcoBBM9nBn1xuBlasWsMYRisLRc
ZvEBQns6JL+xxyqv8TtNndEKphyDwX07dxHqHHy9tyWvCc6lOziZvu+OWq72eanZloWzMteWFNo9
pfFLHUnG2+WsEj62uGDbEoAbgPTCvPlmXwsEiRxTDcCEKZNcNIgsz+LattQHNko19U4lFgHRlc/r
yTnaRlz7gen9V5BQI8nxVkh+/Mj8y7ryFDl5OGbdA66UxJXxbhR1adaOsMNhIeq0otCPXRAeEgOy
hbnBEemlOdIoWG9vvEwkW2tTipq0gorVmu3KB9scjfblnbXCxJTzM9wf6nK1sGrUZVdYOCYwrWLT
80uLFqJY5NDGIp9TI93qrU6C6+VkAu/GkTJee8tOagLqoLOMbeyLmDt0GmAaEd4AxZdqXIz5gL36
RnzYv86QzbxsxlSfEjQRCdsQ1XJPKjuzQTWwml6r76kclbaXFhpLghpm0OLKh5DhOOkOvDm3rnRN
EYX8a/VdSLS2Ufj6YdbdfK7Q3H25tf8LURLYrJodAL1uoYvPdyHZtK+wKxvQR6U2vQwRW3edY+zv
ngpWwZDwsycRt5Rgh7UXund3DmxKWbxiowwuNsVWgbyc2LztZdlR4+jL4pndz7nH43zVuW5/aBr/
xwGEkT0/qyYh7QjqlenogDe0UL/D3q7Ia1dtGZy6uPWvWvqvx394mN7UClJGWbg1gIOUhNfkPtQs
TiUfbPWD+ZFH3vcUcHuNhD+V4Xlya9oi5kLmt85F+ValSg5Fhvo+xOHFvqbTnYBAXgDPPxi46WyW
3UAiCmPvQt+bMCNBxKxgOMu1YdKgbmdnj5qE51zZwT6P2U+pxPKOwWI96gBKfQ6Du8vN5090NoLB
hgaerYgKOtqGFrZc2SgWV4XWrYTgIaGcGgnP3KKefZ2wXbfwFbMOvLtt39Xer4JRRO0qUrhteLsM
ygW6lh/xFfmB6lseW6ZZsrhQShn7ZhNyAngybYI4/sxZXKb99X5MnZGatR62d3I8KGFsTDyWJ35I
WY/bkc9Z+4T28AntC7KkZqXau+s/3FptSQj5oKmbgqNHGTJ6mf+b9cEAiOP67trL4T7VKEvVf1Ks
qwxqgSLLCpPLe9yDzXgv+t4pVvwM2t99ukajgNBOH6ItksbkhH24EiZkBZsp/+Wl1UGNIEXJfuBS
B+pA8B9UTeOCDxakOtjcAwel1Ps3zKF0BUaTWDR0WHttRe/+a35SLrazSHnu/0ngbSrfFGwHP1h2
8X2R2HAsGkemOcUOdInItFMdqgbLqJ4p0QLh3mtIy1q0d79Sc6i0lZre+kw5q+OROl+TYtKJlgch
nXBpWE30+m1iFCm47G0AuBbo5HQTrbTb6GrJlhn6q7ydDhsH1zaBo+N/QPw3U2vxZ9YlfIK1sP1+
+EFdleWzFR2TwLmM+v9K1H0d7exn6X827RiHvZHlVh1u0FASe/BocuhRf9iaZYXldxlTXociM9U7
Ni67dEl8sdSKMrIvcibhYaJGjf19a9kS6REur7WsbAjVuellfRGLs7k+7lK8AhugWs/YRGOgiT2K
s9lUySC5OBQ/UAvjUKxsFuEgw1iTOtESKzaru94Utf1vQvq1H2V6xcc8kPR9EBOFJ/uKGRB/jgQv
ms80D4dU8c/naD/fK++KbOgL+QjPgQtB4EwlHV0OZGHfprsiolcO5n+7bmZZrvrc7AUx/qyef1t9
y1C2I5+MDRwfmV8uX0EX6pF5AOvNReZrAAvsRxWYyYjlsdTvwZqAD7gY3QGVe9hXEreVu2ypYb19
H174xND3o11H3muZwCLPegYFJ0Ttym8p6QIQbluvCxRdqC67tOApGF0ZzVtQcxkvj8WIybEgVluF
NH0GNqddmPgVdw8M62X90TP7PqAMKXcJVJNTS0iT3B8SXAU6CrgU3D5nx06BMYAME5SsBAFET48x
gQ68fB7VsU+ZZ8CZ3eFuahxZIqqWTGpKngGSRiAvMxiwI28mp3QYDcnKNwmw+8oRqhbEWKTdChVD
CcyXK/600m5kbrKs+zuZRHR4GuuwvxWNkY2k304AyhqoicMXf8UcF2Idil5iIBU6XxZ7mOm5qrGx
DYpA1ULUpC9Edl6JezaX+shitaw1Tw8XTTkARAqY0fRzz8I2vKTGlnrqGjj0Jn5FAET1gEFFb6yK
VmvPOMIIDFjazBcvk7MTzCHCUOohx64VEtohQ6P0w3R0liF2rxMCISY5gxYo5pdam2R94NJ13i9M
io0GPY3aKs2SngijLwtmU5wmd1TNyXxcgeaR+33lzz2aKLXf56mLuX//FtDY9hdY46mHv336s42Y
DA/LDpNJFM4NQ1VtTIOL0nR18HL6+6bG/z0jwVbXNtf9RbD95+h6YH+ydTKp0Lq4KNAeWOgTkmFT
S2sHX01FKCCSnLPmam+uIqhgMFdtRExQK73yimdpDLZawnPNXglaqeObf8kOgxkQJaMFQBNVhFac
1QJSVbKtIQ6Q08v/VzIq+Jf/zuSFvV035YhEFfo0/BXeZkAIt3T7TIkTEnwXpkKKEwu9RC0IiEXL
KRJ2FUIDrZ/NE224Bexa9iTSA1o7lkA9wXCgj6rTXxuq/Y7BeBy/aHUH4DjlCTQhPAbk6s26lWTQ
sZomF3n0Hj4NoUWHPeR31JLd6HRTuu/BftwpC2BOhB7EOV8k2Ha6JULinlMGPVrzPBTlfppqUo90
v2JydOFIgQNjbJvpPYNlzQjZwTHJKN50p6sJpNZiFbIQ/yXF8hzlAy4KbOdV4fTX6wGDDjX+M3E7
bprsVtqUGWvL5FZr7VeLGtyNNCbQrNqd7PePDIEg8Nmv50M781ubIwtDBaAAbDcgPOwXSix0Z77K
rB898yWIp6rI8ZDBUqXTwCaM5vBUDJ1t0rY6yKy7EowqXsqM8MUlp9goX0sBmdwieKqjxVQ360Pf
ij40SMMMFk8r4UweXdak8CUR1pk0N+D3mTm5TjYGz9lTf0r82J25VQmBDjpSKTBtUalZ8BD1LZuC
Sm+YWQeeQyFXBZuog3GtoIzSuwvWzTUJajxvVgbBV8jHTerI1FnivKMMAWhGAGppWg9HfXMN00rK
4VTNa1G3NUcW8zGX1zEvcZRMWohgeZP1jVy9zotn4Jcf0azDDv4Pi8d9PF7Ma32CID/lGKSx3O5M
0lx1q7tiQuSG/xCTLimWfDxZo1XgIPVmohHupLPQTH/pmwl0IsV707uLPdiWmBm/6SPgpwxN3TN1
JOKA+C3vKmPYyZQEL1shAzNqJKenm+V3zRTHl/eKWsIDQ1crjpYmmXB2SXFQk1EqjSPzHHELtBDJ
oI2ZW9qhepWif6NJekAe/oVhFx2S6/Nh3GCa+sc/+dF0SpJRfS3XKAe2csaYUD9aTVAQowZF/T2J
3ySprCW1aSEprGFBn7lVRKOBfKRVlQkPkLzUAJ2l6jNkeTlSodhyygmzbmGvXM+rUsPWr5mtnBp7
ydQKCrW8TT3npKt/1zJ4TCMZs+yS08/mgOC8pOuzBkUih6I0Mx+XSwhZJdnHkx+t1w1RTxLiJtI0
IoKWAqYrgjRUARThcl1gb0tFBfI/YOD9ljqEfJBXmgdkn0MK1dfhBjWAmgGLkO7/fT/apjkQMf5j
ye84ncXhuya8dkKSoK8qlYsDJYS8SCERCjlhiMgT67uKMZFk/dDhrGxU3H7a73XsLOc5rM9ElTnV
OoKimK2Gmf3sZZ1SDhi9bWiXS8zRfBGX2xLr09jFi1B2lZfFO6/Z1ssOKZ0Gvx9J9att1W//Whhj
5l/VOoP/mn8pO05liWX8xoFSv/SSANSSfl2NCh1CKXorqF0+SADY+23L8YrRTLkUAQ+mcxzx3wU5
ZSrt+dWYAswHtvL/cVOQpDDIVTRcjYHH2sB7SLNAVbqdVYk9B7trZ2CpLuYZO05Z7Ldo5OkPv0+Q
hibo/TuosXEYVcchEg/NLXWO9IsvxCrjVx6nt+wA2mDM5J7qIFJNO1hHSGUpnmN1qC6OBfmEUm2S
0wQPRMxLCISIg61yLxa8H4yLhkw7PowWfzCA5Nmy8TPvG2REhTJ6nC/ISjfSWn3/NhbaiE+/GM64
mLceEmXslHKhlknEXSc+egpbq0UVuaoyQcnuE23vzzMk0U68Wee30oCpaaHg5NbXWIrEpiGEAlVS
g44L/8j6GLq60QCuagrn66Gq6fJofYCczQRYFK2esg7kohh06LbW+m24YNpKsK+sksSrB47pARxa
pZaLCLSnrs6YGNmvumN0dohtmmRPwjYk6qyazT1be8udGM2Vl1C3gQrPtSKJuzdZBnFmsSQwd76d
C2xU6DBG0em0HvDoCayX/TIIH5LaTCwBwhE7qPS+2TJKOVw3NrdcLZyxveb5bWPMXaOdgwq/ltFz
1T7h5ZFVp4DGXlm6vjgQcOSEzweu8xuLdzhZIzhYq6l9qwsvr68H4wAEzzowh9T0nBy2Bx0f48EB
cURQWMo4lfMZ4KfexppO8KN4d5JIWpyQSxahaLT4C8SWp0YW/1iMiVBrCzQJtlQqDvowGk2Vqcn1
b7fYfaBfIrNLbYJWVrH/5hYgxfanLARZpDaK/Hu7wsxZtbSVb486+dB4B5jdtU2KrUrg9hBz/0tb
w1CD+LdK2eH2hbJidkj3kYWaavu2EM+LgQzjfCMi3yVBruPEet4znxpu1abdPemToAmNbRxIkNsT
31OvCWeowQ1IksyyW/sA3eQqgsW6M3xsYyuVk/KmlllBX/9fJqKA8588EuNUNSDfOhbr4CToknyX
lqhgAyCN0QGucHhKd2gStkHw94QX9Ja7XQQzCuXSg1uPOn7ovtR42g0CSTyIQoZXidAZHZQxH/mG
Oh16gYAgstInYJAvePINdIZHLNJxPWOK4r9NMBKSklq9+fu/8fFExZ5w9NnEpYTEIzWz5G9S9F6Q
PXUUJ9uMfPCb3QKsgp1/4ckxBxoQm/XlSG4q0K5V7+JHtqaqqBjHKkTbEYC7hVU+Dwxs970QtId/
2pdsHXPRI2ZaCINPPBAM13aD72ZZBo7a22A+sPlQfxM9w1g9oYlhFtO1Fn+CU+F3nhUD1u3JdxvR
5ulYxK0qScKC6MyPJQGABrtB8f9SEL5seezdn/780eQbgRcDNB7eGLWKrQR7XEcHG6Hwj+jYFhoY
b58Q3Ti4dv4htDkoklgWp2K2G3AaHA+JWdHMCWxSqla4qvHrNQ4rs/JpGtpsptsFLlaxH0RRZf87
yMkc8qW2jEL+VrQ6XKnF7aYxPTHwIS5LPlXr3JKEcJMnt1dRUAIhIrW413CTrOTf9Y7LUQKm41Sy
t40TuPjmFOgUqyPxxz/AuoNp7pbTkqDwJpWeBM6h4FiQIZel9iiurmfZITvYdXpsl0lj46qrMKpH
UBs2xbDFL3yQ6U6MNR3M74StcxrnyiQm0BdVoUTwRtU2GWgxfuTrnTmcQZ7vphh7zm2JHPT/mvnT
o0ilXF0ZSmIjo2lE4qFVk6qp6lTQd8DaPqfQ3nWyjJe2xYdxZa4g4rUFj7dtq6q6w+QbQVhLcfEL
lJ4KOVGDdcy/dC01O5Qr/zYfVtbyThJnZB4QBb1OTXuRHNRCk7coLdnpUhuCHq+LCS2m8kxIqa+i
7rYNkii97TrT3oaWu4f+I7D7nRcHPwI0ARO+4lQQFTaquZp1sMe7l+GfVzm/ZPk+WjVw81DUBxAo
8/kM8YW6ZYhcYH2+CXqOKRs90h8FlqHP49btHI1blrDPpjIchkYDpQc4pKA8+2KSy+tTDOiP0new
nWdEFa3cEHvFgylRWdg8zUa47OiGediS7lAix18IRTC6DDRr5XLvYLpCYrTHM7VrDb5zTCKsYiuu
NytEcwTgvnHVH8VsBQggwK3txv43zCahvqLmyuvourslVGdW37AOkiD+jwKXpNlhaPRF/bq2iVDR
Au2o4oaPQBJkJSzNIAEsNpjiVbfhIg193caGcp6oQpeN4imu0dxJOeHlAYCaauwsQ+u1burkvxNI
T1TB4oCPKraI998AEyaPuMwUi0wJhsiNa+7LykC0uNnRY2akNRWn702xOHxKl/p4qhGYv2brKz3V
yptOeH4zw3L/mRs1wx08rC3FJkXn0S9gxtyb2LAsXlA0yXGneCDjVRmxXAdLAGSeJywonzSGrxpu
lT0Vfwl8SYMvCkOeLUVXJovtovEw1wRUBvk2ahNhSyg77RqXAv7omJgxO/zfZS1nEDXMYOPan3Ui
2ch/uPYDvP5MIuZ0eoUa8i66eiFEOLhNHCilYyBtlB/MZSwdzLNrId3s48HIfNEQd2p5JXqqj359
3tX08CSjTONj0EgzuxYTh0iGhETh9VuKe5/jhT0o3nmF8xzFNM5/DccOhgcHbE+mNt4Y5U9hweZx
DnbjFtv2KuLMoG1v79bMXfTXcdoYsdie5jtZ98scbT/8piMRBcHnfvEXZs3n974SsUKMliTITC4L
y2RYT8MINJpOtHAvc46+Vry2wd1m+qbJ3AbLb1FwvN6s57TVL5+seXlcjXu6bXrQMBbMWH09KsDp
tV1dURXpxuWXaeRAMxdN+qZZUlE7wREFRy44KsncqK5iLM4qn/0w6kVzaGWj0gRrrNpkINTEYdOy
0PziYOweIi9bNic0atjXER+VcswIbLelxB3uttJPPKM+lIFXDGk6yuUHQ7XgQ/OnKwGoZZRLLXLJ
zU0L+43bevo4FlVWvSYN8z2ks8xdIPtjzguagh5Sb8zm0mcjGAg5PFxgphCoozbARDCKqg47oWes
tEd5JSKr0aDMu3gCDi+oPozkQ2C22sIiSP0e6dXdyQsYCT+EXbj8yMH+uh8ADio/Xjn4zmtUs6aD
XpaKO0amn76s/72nf/9sYCOLcOHeuN9pqHlw3L0Fwea42CWttSpZsKUoHgRYPvmfge0jR9FW1b+w
lmVtJx1Z1Ts7sMcysmFTNZ8lok04GGID4CnS71vNZNgA5SLds5+XyyR42tiEiXKcmjXPLEqzA1sg
cqCixOTvB4FOCmMgbGk4XnqIyf/4sv3Vm5hCWqIjOEUCxeVDZUWep6SXx1y620TOxUzRVAdzv98e
5u5RFbVPx+asPAvxsanwcKWpqCb4ZxXjif0goYwiMbyj9iVuHRj0K6mJd87X6HOIwRapH9Ly0pYI
g1+8lKgV8/P/UA0Duzq9zGhgRBpsZ7kPTHLfydzpFcQI8lZLATpOJIHuXQM94Sm/C+evwZoUYvaZ
riMXTjVFnzUWmZ9NGx4HgoLDMxu8xeejZg/FXImfgELF1DMwE/hTADBhiHki6lUdBh4jXr4M6Mo5
zWJgBZw/igsdWHAYqdiYXRnHcyp7eh4vaP7cDTX+A5rnHdFF0gzS0IUUlgguU8SF8BFC7RA0XdKb
FU2VARBk5L6TSeqpg6CJejzt9utoZCw0xm5bKu9/LaYcO1UHLJ5yeNFUk+Ds0Stpr4OOI0P4/ZpX
3IdZsKyShYRy9YMQIzz3MLTuGc8psKEcqobo6jEr59auiHz5ZLGImbsMHWY04hoIgmSf7OKUI0GI
Fjf8QvgVsCRTxLxyqazM9+m4QBjmYH++zcsT07a93KqqE8p2m70ZF1XT/dppzeVAdjZwaOCJmDUW
X+7hDEkBkJHUK02Yr0u8LgGYBNUpXw0XQNuCd+DQAxgnEXXLBjzPqXujJRD/lBFK9JD81wXfNCYQ
pZp2fE/DyVH8NVQacCm5tSUncKkC4+j3PAt8y489EQQAmfnKTy4mP/lmPJGIjWCogXhtbHU6itEY
u3P5CgIKNkcGhpMvNo0HH7isE/4/+1MCnidwrL6zDrz/mmXU1PPsMvj3ji4LfRSBUIDnngxPyyH+
esEbyrFCrYTTH1YoXrIzqSQ5sIR9di7rxyUQI11/i4r2EEyHhA9JVn5jn1xjD4z+pYKjqBkIN6qA
9d2Pzu17pqVPQCEH9DG0mURAy+71yNPkbEFntQRjgfVsuwRtU/bTvpDvc4kpXEkvX8+rSW0cswcL
OKa+Osrg8zAjB6b13vlpXzFGIl+KR9qSw15wqKeP7rBsffv9MXLHNOYE6FrNi1qNjcq9u+/bKiWY
RmF04Y4BtP9MpkcU4ohgo6Yqc9i49DUSU8lnX1y6vdl0YCzI1eSY2pB0t5Ygqw2m4K7b6QGTGDKz
POYBzWSIF99jbZRaxpOTO4nzcLJtxQtFc/44p/gUr/JbleB3zFUxKVUAxFqXM5mo2pw50ae4ZMBM
Wyoh4nr36F9Uctr16Amq01u/V8opFGdNag9pxLu27oPsV0UwkR2anFkorndlo+KKmBCMAh1Vvs18
5Ys6TVN7uCowl+Q0pMPPpJ7hwGVoWLRE+AF84nIEEHTM42P8w9iF9fve20Hrd9JuM13GKJAI2m+Q
0/HhLz/b1x8znWzQi8DUCdT1lnF+TZDCLqBZ9Lxl42esLXB87NJn/njYRdAR30S9wUj8LIUAjCLW
RUKQQFL28xxwhZI2LnXBYMlIEHo53NljpZdaPI3XICUCEs9yN2QLQ/3BWFXvL6RJmdCbjrI9Xy0m
ILmLnjZUhbHkMpwI3Nb9aFAG9ehi2JKpG9hZGlV6N2afmMRvD6yGQfd07KOIKhgUkek5bNdFgSSB
MnpsM5RAQ1WP3t22rqcxbPMFDkuCI3ldpXreNcjcxXHeCokWVbb2mXsEJSnxMbHplyotSIGqohu9
2N9idJvNEi1OaAkuQmM4SmT5rN+knL9qAP1u7yhYPwYC7ExBv3l692sTBd5e/kUUDvRj8ua4FE0/
hTJlPdfFY5AhLxP4i9pj2EfyRKRGD4cRK9yuR/5A7ffuvPTumI6oRt/PUcYp1IUnYw6xUVSHVn8S
9GTLm+VjF/zMjQPko32WL07DmKqCjtxYjLU0kN2SFh8C8BdimjoxuahFd/TBPyNbQz2rKdpQ0Jsa
AtrmvlHGUpgNHphY2fSONdUieZ7FqktlhSGU0lBcZaes186QOfZGI2GHXN5Pa+/UsZ4kca4IhMGr
f3cWYzQqcT7v4awYeAkmqTyf2QeziT+dbGkU3CbmS8mYDuZ7ZqDg4K/8HFMt0oS060h5q3bLyQgW
x1j1FFrjBDV6XvpO0xFEbbJhx3BBNfzuSXg0dg5reiHEccgFshHu/REgkxiS5rKKDBmnKZmDG2zQ
SmuueLMJLf2YxKonGZCu4QoCvi1RRoP1+2/r7JUsJdFExySRkY2qzg3SwT5fAklau1uJJMmCQGbM
MtgW6TFKL6RzJQS8qzBxkCkl68wTYJQQDbJuH7A/GaikuNrARvaI4Ga+oYWd8vEjErOQryt+OYPy
+zvljg/NifrQNWU4AAC8qR90N0taRs7PZyQBLxZataO7h5v6u3A466YdIQoJI0PrKwdPOvm8KHce
NIwdTzyOJulZQDTA2HaJvvF9klG0+jsaBqTM1/eQAw7jw1OKxNYxC/38lA4mJiFOn6MAKFqU0Sxz
g2xDjzDh0jwClWRRUlQo0gNNp4J/tgsQOyhkPnCrsU/syuGYgr54TRDb3MCs/TWIeV++Wydol1zO
/TlHvP0hVWOvrLO91Tq7uX+RMhv6Tn/BhCHKNgKKeO/OK0Gv12veFuIzzcmYNAwf2umaUtDi05Va
MG0HdxFF/WcK2/ypL5i4ydW0fFMbNGrdEiRzNzWr9iF6/vH9SRMYTunQJe30Xf5CMjjsCkhXfKcC
R30X3kOIiL+X1yQ5uUGCkl7/kokc/1OiDjQKkdSExRYBasg9k7NXZqSXFwNBgPN7Kz1ypk+0TJQo
sV/23JKLSGPv9WFvxByV3Px14nuFYnuOPnQWJKUkIwHzrUWdxf4zIrG0IQRjNg43CcQFMuqZX+Cx
bnTxuADlgL+QxVMFVdeq8co1vqtDknsFFMQwro3CG/lVSr/L7iOnJwjNElECbGIUUyIsFErqXJM/
+PzZNxl5wpYVtna9c3NqW3g47sCsU1eEND3GWb2aVImOOwFaEZDAITMNBzPwvXz/QFZtR3MLNE0q
bhWW9EDYzYxrqqVHVI9V3ZRpASqDKssM2TH7whXoOZsb5MWq8HznTqYeKfNQtwLHOZ5hoVgjUolk
bOYjAMawNVIlgXKhEbHPzGCM540tHUdqLJDX8MZpw6g51jOyqiW2+uBUIe9O4AtfA8TZ3TKK3m/2
aMyQe37MasBbf1IO+dI15Hy5a5ssh7UFxs6nRHhWbet+Q00tcF+MoWfqG4aCj2Khpom3YBCgNDtI
jkgRioF2zTTdI67eWBS7c1A5OQmPZT+tgc7VwJ2fhtbVGat+ZkHpalNpDU+6gnLfAYcU7k9Ju2xS
hd8xLzVqHjgvIQqG84gbrUOuLH8ZqBCbKok/j8/4oSNT2NJOtlougSsawiIOmkUIQqa1g555MPG7
bud4UVIfRi7Stel421nsY2Oo1Zwz2cLVHWck88XbO/mzsgUzfn3VNQChohVfHXAFOul+D/iYFi7B
Ko11LE6Kee+w/Wiy8oAq9cfrYKCaWEmHd+iPDBLoBAYZOPTT/neFD7fj6a6PUJblF3/SmaHZWJwK
CrhekVoYWOUpnXFOOieuJRlLkr+FkQZ6cLYXkBRBoaHBtQHy4DXOrp/pNpILCxowsttJMeqazKRM
qtpVPT9O/f6+gE6DsOZUAew8GfRcVASLqfBjaDju1UiA1V+gguyrTRK2vaYmN2AXuCJeOKuG7ls7
syrxjSrnbEywaBWtbyzU8Oe/EcFc2TIiRm2Fjm60MhP3Dpo0iy09N8KdSiC7sQDEHqqGVFURQwh9
mzVSWtOl5U0nSqCBEkZTEadwicWE6Z6DS9K14hnUakm0mAzZpSAhh6H4GvnMazRlkkRFe50JWXJl
eiIGt+5dF5dTboCwcnyNSBMv8fRgRNefmux1RmWHztcl/MlnUt0TE1uqDph1W64IFbrkwmy1Vfhb
Az01picojtrtcildAqxBogU3rxcmU9Rdi/w7688X9a07vMoaXEoMQ+Z2/rxaCFTcI5+rvxiChIVh
mTobmxzdBGKwpvwvgIBq/9TAsdhPxX3zHmsrHYgu+ESnSqEJf62BY2fOWEsnTuATm4QpsPGGFgiH
T2rOPkyIaoHy8UREpwYO10hCY/rpupPLcZ0/XcDW1v0TZWh7L+9DwYRRlBpu44kjmYgo2jVN8Zfz
2DYKFbR1SZ1E/uibRl4yTky5SzEcTCcVbvBvmqdjhwPGIzoR/kL1xl8EEFmliNdmexzl/TQvDjsb
aO7v9MmVmR+lBmboM50sMFRrPjbp73UyNQC1vg72NXpzPSCwBwowNGPbk3UGvIxlATeLuczQWRf+
g3DNiUie1WsA9c7sl/b82KhG3wnCI9kNxU4GsRHWogkgASvMUx2VfF9JfZlbunzk+/iZpxqHZsyZ
/HM4arqF5HpU9/xXNu+pUsJJj3HUjpIUbdWd3/MdBNgadDTozOgfZNM+L8TuSdZ2oG6vHK8MpsGV
oY7HNOwXxtPHjZI9dRBMqwpguRowcs9SOK9XpbMTYQYbFTRF3/Yk+aVuomi5nZV+3mil4Upau7+i
ttmIGt0rnHlIurNXSJDBhA5pMseYKNRriMAwYFd2wa/sSdCWVoBceV2Fxdvi0bn9c3q4Un8oea7L
VAtUyn1IJvMuQQaOhorv54pZBgdESfnKiby9IsV8p66BS71n3zqFwHrt8lkVtdp9Q1vBKr7wrZw4
258PXO2kXNUoT0BnF54BZOeAf21fY9mNtzAeRKkT7jLGq78INuYzoH/4FluMAgQCIOyL4fp7YeKJ
8NemdFnJiuopJdIStSstm9KFA854bPFMq64yRfxXZcVGXqEWgsfdAMCVfcpVvCMf47cYkPHIGky9
dmFwSOEESqSs1ytR5ow2ZKbb4yTRgrg65agYc+pNP4ExPEUb9r69dUJO7FRMr5ix8iTGz8hgVYNc
xbaCLJZy+26bjW8uJrM3ODI6JPvxrYH1sxe+V0f9DQYdh5GZbxFVEIatRVAtJwlWc775aUgZeI/T
OpTYRJahOVEKfCIzk1hXlN7m0GaDpQqFZKTi0syUUnDDUu/VVxgYml21kBvR1O5PPXRFNdooNoAt
yhBQ5jpr/vniM7KUjXb97CycvhgQjEaa49HPBg84Mff5/0eZcaqFLiXLqjHzA40S63FV8J0wtD/l
nXWd4gwOaIwzrZZJCZyQOTUJiP1FbfX0c8416KEyTVCBByLWF4+1YfmGaUzU1zc/H0meexIRzICO
Ma0hBqBBEKa+3Vd3HrDu/fUWzhb8MfpvOjujQu3A6F3VNAkMWI28xFCVVNc7zRt6vHdn2lndOFkL
e3cfSfE2WuBl5IARjB/nRZfVHPhw1gtJAI5+zcsx9jtXsSGhVkQBIFl9+GzMjSGGbh1pBs9od19H
IyrEpBRIPeMk14ou6g4zq981aIwMcTuJshM4sSbJdtfWQZF0m93qFwtgQFweLuOpSpW6sxBOL69Y
LhqhMLiT92u03SVVBb7PjNqDjutSqUifvO9TDT7eT2utiwGEP1THVXBJ0nN24HS1yIMT46fhkaaa
IemI0BIebvW9lMIU04iwXXjvukurBhsUvKi1inQ/MtlTsnO8G+wtHCH4v2pkF4XOIfgQZxt3w3Xm
4yh0u8Tgct0CGC8HD/8Zl6QljoXsLI2usqsSboO/BKIpHftG3KSdzaCwiZls/oZENZFOHBeVbQHt
ZzIHOX4Q/aqRF9sJapJM+kQBjT3ofTwsz800OVhcWY7eRVIcA2AVmsUN17lbBLeR707yvT2so7cp
gGw49qD2Wjty172T+09lZmqb67BfTOtGbR/IYrIlfFlZfbUSP9OdDFa4gInUwMuxQPgy12Kn8Be1
/UvvwvhOvNT5FQkyy6XrIX+q4lGfJOK07Mk9Nod/SjCL+9qaP59har+XH//B0aPO8n1toWBH7MHT
ron/0Sugeb+l1Hlh12UscvFFDaCCUVgssAmVDD7aSzXZz7JSN3ETbAkhGDcx3LXDtVTo2z3y006C
0zW5el093NMiDh9Nlz9YxBCSIyMSoy1ZnLUCNTvVkg71jTY06NwcP3tcJGPgv3csdBGpE0L7Vj+r
GK5TlbYXlMtXueogkHKruYRFt9Uz0XFAVSAVSJKGiKkZX6PEWd0DIU/HPNvEMRebdwkYZqPadu1x
VTc7IMeHbIF/wTPCN0Bzk1Bi+abdwEsGkpcyKArCLg1uVuwKpGOiDzvfPKGnrWQrDHND5gFtpaWZ
ObGUGTa64CU98w/sqLmynL8O0nHy1cEt4DAgDMQaHQidaq4tbFGBI78GtEsmvzaYcBR330MfYd4m
2qRbP+7bQgU3c/NAEwXbsiOnUeRAG6HhtDrdRaEV7YFu+fHFj/EFrr+HIA7m3A0JtZOiIJDMRVyS
BZcPtf7uR5dOCLg8RdBoUNjaRf11jT5Cqi9u0n1gMQbhoNitxbe6iZD03QhydubR3COu2MO2w8bd
jemRzPz4vyaY0xcHh7pAJihZ3YyWQcybCzaiUx7wMQDzABf+kioaTExxeFx191Rs/ZfIakTiXKAh
Qv48OjINi5MYNu0o/DehqdY2uN9HrBJ0k6Xy7gYNMeR78jYNeWSHDc6i2fI4HAh+zF3ZsXTtt29h
R+7DD9wtOfEJuzumVsrumTCOGLlJBWbczUzK3uEJ3ZXZsnDflAwx6nyRRT0AZPVXEfLDm/yWPwqY
D1iF8YCx4tl3lWu2sbzdBKuxCXRidAz13Jw/hgqWgLmEH1+q+t94vbepavGSFlg+gPg+IgAnww0e
spSsd3GUdtsypKZWJ0ZTQrZjJU5u71q6PNqSFk6uZop9/3IHfPiqazfbQSjmJxuDoU4dmXkgbTi9
f6SjbOjuFkmMvh53tqed7uDfzKoTmerepXskZLuDNz2L118CvPJdJGMR3YE6qP+hN/H5nZREjIS1
B4PARaD6uQs5MgBTBAlbpxSDPkmKJWm9tPgpaEUDD9U42Fo55XJMIixQfOXNsDSGoL7w44Ma3BbZ
7D6ZJ5tQ4X94CJ7CQi6tq9ZQZU3C2jPw9WjPSzVZpb/GHwT6MAJ2lIIACqJp2Qbxd12E6Shgttj5
fL1z9M+atyQXfbXJdkP45xlFGVFrsDDQaE6HH/81u9RwPOwdYI992Z+JUW3NLoA7JVwMAYpgkk1X
rTF8/Jc7fJ/id5GVUJDJiyrbHmLSpuuGGpasOiuABPyEQFrCxd04jgSBpe8YisqEEVpivHgZDvOS
NsAKROgUtnGxHDmZ4Vrslbs0ccyC7fLgBAwEVHr/agN9EbnNV+myC231FDNsbr5Wm8k4awpADniT
+gbA8aZVYAFblm/jiLSOdACe0ZjuAFwEJjhogUI2ZEhl3a9RNrn57Djt83XeJrMcvxP6vR06rE8y
gG2HB0iK3ZqE3D6AflqxLejh0nDxbiJKm6YMYf745nb4g0P0bK3Jup+EitVhEw6zhQ7GmOBz1b6y
vu5zAij2aL52Q2+q5Dt5I0CZLwCayqL/pEdGNo+Uqys1pL9PBSITnwRcGD9cU5K3Vh3kWYhtkcIH
i+7m3HuXnLSj0o3R1EcmxXnjqFVN60QoruUaN9ADwWerHt+Hgajqdx201/qQArKtmPjoB3vMfKNp
haSpSZbYzmd6MCgstDpE7g9c9YwP9S6pXen31vUCLO1y54EFauhXtfknWGZXYjMhXKd+zjclFfuf
lI8lbXxsoK85NfJUP/yx0YNurlI3aOrMraW1RAeeDWrOUTw/zaW6d87JM+FIMCqaUTvjymMFRgwK
3lhaoKWLl+KxAZj/3zVB52y1NhfUmnxN4fgj+8Rmh9ureaoWlppZh8UhPQP01LqvMv/0sPylZyIb
r2D8li2iDWcPoLLAj9F+S9RoBAVHPYbIsuabYNf/m3YgoxxylpRb8hImEaLUWIqicxiOxOmWZsXq
okX26y5GR7xnrKYGRdzf5x87wiHG2O2R2eIkW4aUmPiZXW+utO8iayO+3i/bjICjRbJkpCimkvlA
wktSP9lKdR0RzMJUXhtbzQUCFSfY6XuODpnsxfzocTlSEQSjSJLajPovj5Tussj1GMJCh/Qzc4LC
aktg974dQOFjxHtwlXJvwc2it6Ll1XLouv/5u/BJ7xhpB/eF/dSTYmfOChoNRGwdCRtu+t8EZOQt
bIkcn93S9NbUmm8mv3DPoiT5HGF+dKiVTaiDf5s49CsNjCjjSMdhvHB/RVdOwohRP7dGBJpK3NK2
t/fVCoD3qPWHznDIIxK2bXbXtTXPKGU4k0TZs0+n5F8b1BYGA7STkn312sar0iixA6z7LudAhHwZ
cMIsug5+FnqZ7QcUoirfWj6lQIEL38VeZwIAzIoHap/JtLco7fqdT5zzuyKcXnHtEaqr3wIQHee3
7amQmZDAX79zA7D51tfg4Queb28ww7d6L6A3nqjmT0esFz7ThruFJF4jX7A2kuqoDZhWjTodUzQu
ZcnfH4UUOOpmzB4LsXaqbyrmKbPJUXeGJF4heElLmYnjVyex3GM8E5zksG52/9yahpcMiTFnUhPs
u1JdlUB4CfHQrFOi0vvHcu0Qx1V9FSOlq/sjLtQ+5MCjGfW9N7mJVF5N+jHZL5U+VwWlKkzpqMCG
94V8WKFyWy6uwGQex7Xb3Nltf7d01wHpUlU1D3tGEoDQzhfMrUKQyub+NoEa/QOivy0vRekw7lDj
cX42Hs1++K6dWKHCqdJpLqwQFEL42CxY3wlH+CLi5Fm+VZHtwN4cQWGu+M/WOzrNXJcAnsupZvoU
Qd/JcEMbxBxONH+H1yZRh5fbdAi7tTzn6UjIxthW26lPociytlnKUuOfzPO0uKu1mXcfOCmIg3xt
fd7W2NwDFrrxelLPXMgAZBaebPGhSUQzFDhsXPbhA8Jg626AlKf1/iNFTWryRTpv7NeJhEUByvsI
Z7Z8ni78pAzgQgsOMTK/1A+PchphlT8YABuwuOnXn0tKH5WiBmgE4VgTCcEsWZn3cUV7OZHKGxLC
+ZNXRG3eHdGNt0aWmDyHF22X+qt8vHVxOpHhEGeLKlLnbFVu2k8wqjasyGFUpuatftjpAMgbc2w7
HVtfVjxqORVLR9FByLKDhY1u606f/yfo1slJ4n/37ENnF9z9Sz9zyIKrjJMrdh7oZF32ncrUusvx
7I7wEGjQ4yHDQXWDtPhGS9GcRSeaVOC6DhItxTqwB2O10bHiGQjdOPvsU31LNxhEllCxAx3sxEv8
pGrqNwkWqRL11XR0zpri9nbkQMhnW4Dpw6nwbS6EosCdGSptWbFb2WvXJUkQ+b2j7BL67c1pHNp0
Y5aeFRBE2CU1E60cLTNxzQJkeIs0NGLaSGwdB9ROYd1HmSeYhrZpbb3Z8aC7ho0ug87OF/WMrmby
kwEbgVg8pAmNQ1s4lYo+YGw7d8V9IlHOKwdqPAT0CF0tr1K3PO+CmTrx63JHj2fNN/iDBookZ198
y9bOaKqCBcnV+1ETjCj5HOU2epUGcYgeOsGnS00a40FQ8B5MOaTC0CGoaX+nuEIl54rYH9ZIQKfA
4Mxf1RevT7atV0m6MN78tHqenDmSBDzC789JbrPShEMNzqfND55kP6jk6xNqu+jVchnjoWOcmYx4
cqnX3rZKuL+keoSWS3058owbbEgoTCJzuQscjqgTFHEDvhp/hCknTHTMaD81zOqJNn1fK9cGwCvA
wFMU2Qa8Wfbh8e2g1w3ItmfK6rIZK+4bxa0EfFavmTza7ZWgfi8Sbpoe3HEU+C0zATKOStESHWFk
W03qimqjtzGdHRha4gZ7f/mX4FrxyBFQ0nzUjsPA33QvsLOYteIeac0QwOrnZCrNYYVXiQSJUPof
5ITdtAjP5nfX5fyAhvqhy27ZceCFK9l8zDh5ynKtqPnskvmkhbf9cdbcwcXfI2fXghFq7GbWCKs8
Cb2h5Dfplppz0/1FTcmqU8RLGuZLI3m7rGKA2SjW0uOZ1sqAqhujplr3NKSQ62zqi5/67XxkzpUT
qVZmm3AnNCj29u9OEj+Xg7wRI3BABZq6sG8qVDxltCsfH7VsAgt5s6UXWfPWXBP1fUaYlZZCFF7c
3K324CzZjvKBCbvioymSz1uLm24DRSJnQOxuhwqlM9KUo5giB2sWuAHFmANv1I4n5sMZNUM+oJ/r
EFCqySqgnGpHVG20ZcUDk2o8bY2d2GcyHqFTPGJMyVl0rObBuq6PUZEkkyZMac/+JfqehUfjJsku
Y2nLRejVtyCdcdjucRafAv6+MX9RRxcT1UVFbOMOZHUQ7fBQ7Zi58jYpYBDOgyvQjQOSa9Q92Rwc
ToilnuF5D187zeZB2U0d307oCadaobDAfdBudR43VXkNPzYBUMYZETfFpSziztFsrx4r1pY6zAnA
ggvZvpRVhM3SDl4g5tAmC6KGWT2acO7LhVhEFDTAsP4ibyHM0NiXk+Hj8drmFNQfdVFzMzgR+SZu
K9GeKB4XZ0cq93Q0XdADizSqUGH/8Sfu5A8RVznk3fQcmHKqxrO0F9Ge9S9vwR82Y6oZisRwh0QK
LWbS5ctWEbrINaLQltXXwFZA2zGPe41gVN8N0TblkhRGjXSVFSQ3BGxeqGvA4Ce/zDP+OlFI5rwK
VQcHjoYo56h3xO6/FYyaZynR5ClAMJzhReHAbEWq8ff5BZj8AwnvPqAHL+PJJ1x5Fo3oh+GFt0nB
rpRgcaFQDtezPhdnUYogGYnp5HcYxUk+9Qkd3tCBPhosPJ0uvCKClI/yfdTQ2Qc6xf13dGTNw4hz
3/+VrFEEjMEbreuc0iN4NRtwAnXRTushH6qOjvVgTWmPE3KlNIHFOSKXRRiLNN0pXJT9FB3026qT
kxNlyBT4x/0zW9nZqytWvg6zshxL+ucU89Hld1v9u1D3CUVDr5kwET819kq0ADUW5PvuyjwYUqoV
wPw08daq+FaE8oXDDAtHO2ZcQvXuDou1lnWRe5Uyh4Mca7O8ztdVXBWFIo0D/5QhT+ACITcDaubI
FK7utqd9ULpjX1H2M+lX7AMYh74tbhLhS774yxmP+vWmBo3pHtdNaF1OPNJgbzrgkcxYDcP66+P3
fbmp8A9j5OTcGHoGDMEC4/kXzktxOd4L0czqFe/SgNvPiaUrcGsrhXiRwqc8+4ysOShaGKHXpG0b
lQ1MoXxfUq3XWNsnoh7Oyvpwf7b3qMYEu5v0Mni4tl+rSIpHxxkPdRCKH2ByZhmrCMR3R1fOb0tT
kcmchs7wPf6VCR9wbGwd+RK2C39xBNQhehYKg2GAMGG4O/xUzbgJozBolX482MGb20w+C6Nic581
q/qHhjzV7dKqWY7PTDUOK0hMd9c8Ni9aijuMeLM1w53OX0qSrfj8KhZwmWveFMvJ93sn/Xk3GyDZ
NI9Jy0r9Xc9CFoIUO+ZsysfG9vg+/n3lJQGQDx1XukXgV29UojBBQ0MezDgksm8Z640P4Cp61fqb
eTwDfwsxhclLTZvhQMEuFbmbTEv17MvD3xW3aWfZzbLJfmKTd2UNGP8NwPuZq64azEg4xBcdX0i6
by7qM1ArRO3IDm8lKZ4wB6sZItjh+vobk2cioIwqLA2WNGYegHX9Z08WMoATEaOsjVZsLXzAm2Ta
OjTqKQbUKvUlLHI0E34215TIhE8wIASp5xKRjbK6v6pNr6t4THgm+4OLVXuvTIgwrnhcWPO/Vi28
OTnaqmI8ovS8NVaZ6F43a2nwZyLw58bU0bIexfHIvMtpoUHPGR+LXfEmHxHqlk6SThdoc+RvxSjo
hR1y2XMP+qjUX0IGPSZNW3vRio4/cU9CriJfB2f+69ct0LcwkU21sK7/v3kLdZx2TVTeCgcNZfBL
plejUlfgPoJMWBo7JQHIpmVD71G//03kBi6QsdEK1X07epL0IT6vH5428tdS5OJwrJtdPlaksxUh
l/bcOa4NPV5x2H0xILZeqXm2vyYtaBD1yZ4L/2C2jEVCwHh/OaM2H1GyRPJ95IUoHBKHjqtQvCLw
Bj7AC6pO0tRyK5Ix9HxF4hhcena+ko2D1ce8eHp1uH/8KQTLxz+Eiggdaca8MeTYN9jXQCdhsGSG
7FT5Iu8ixNZ+N78VdPBY347FCtaBpdElIQF6KlY3RIIeMLbkF2mZS5E4LIuRho9USDdcwqBNFwAP
74vyuflOK9Te9AQuXln3bGw3sX9CDg85MqXpls9lsaWC1YJAGwKkekU/RHv1pFwwBLh22VT25rf1
cmn3ceC+n/K46kBhcAa2SHNe0/50kPHnraFWTl4XcF5/wXczyA1nbN+0bVI+qVlVj0QYm2xSUjiS
BwaKBJlj0dtKy1MWNsrRZs/TO/dJ0PDmX2TN1HwBx67yRU4eRKnLdj4eTK/ou5kBWmlF0F4IAoh3
t/Xqk04szNN21SP9d2KA1JePG4vaFirLaclQLFxi+D8qHvZRF+y90lnTMw5gOYY+RczMRYtGQHsX
5CF396EQg0vI33hMjSfiEoRrS4FwBi3GxtZ2lW39l/3teG4y303vOPXHZafFaeNXNH85Sszbtrz0
yYW+zm67alTbZz+mfjuGNRo09xEKEash6hoDdg+hLrwQfAmSUSfTn98hqDzgzI4/GQ2GMPIWE4PG
kldyTOMvK6TtLFCKqEVPWZKYT6FE/bEWkrSuajMHdSYCtT9RcHIp8avqA1vDwIEhVLF8D1i/77Dl
HM///yrWPgaDEVel3maJrsw/hPt88kZYUlzp+ZNv+CNnlgqYjLXEiHGu4mIFyRolB27DCktwiuRT
5g+jb7usQ1cgv2bmo7nRGSgTtSa9U9sXdsikZkepS+sNQKgvZMqlQgYfTolRHQkXZLOLchwVpgEq
Bj659+622YjrqAPLbaeRlX7gncNOBR5oz77CwmDuhXdjnfBkcoND8Iti66r0grUNIJbO405tdB47
7Il8xvdgRxrPDm7nQxCwWsexHdMxqRYXDQ2bmbhwxMdMtGNg+Hp/AwTOmBo2Bv58PWl4DtKi/e5a
SREV0ytumD5WfzRYvbSc2Ui++Ym4kECJUZxmHmGp8KXLago91oiYGVeAAX3RUHfvc4mlhSy2Mbuz
aPMDrzYBIoDKrfkz3Nisw/oHv6MD319EUEfQvmXqln7Z2+8cA9zipEADxhA/hDbnWj83HD/68/05
HZ46s0AHjWRW6vfqdj8OE5rpmUbDaqqacdyp9ktUXl/TulezI/AWcyQ4xEKA+ic3w2rWNp39w0jY
gh/IgGs5B8WodAS+ZOmDuUuimo0tFsgwEOhbJjLQOXxHQT+1mPDizub5yXY7VFFtWlc43WRZwhF1
mI6N2a1tVvLa8PgXW9kA4ppc3irI4tCwvBdGMkFckIBrIYWE4Gzcu7+p3x4RwvOghRA+URE4fCKQ
GoPUqY/Dv61V+YT4Q0dZ4yWk+ViplB3Hx13YRff2y70n3Pvx3MRnAy6O1VZ8PEbiZ1jgeJYxkggm
LconZ9cyRs/ylW90dTztj2IwKpLupVmffKHjhqUNyRNH/7yHEDgcXAFtgsiRJGX0/EjdMhniA7f8
opbwD3efjfXwUEDVdJX5D12iTlXPXaZITf6J9USnDfr/Nv7o1nMH5MF0i11b+aj/jcCpjyVF1lRd
TEk5Hps1eSn6DdMiKtsrCN6YA6ulhvMR92XIvT6XI/E9MUw1R8U6l32CoiQkkcfvztjpITbDjkRO
0qekwc/4uvankJOhvVBhAqEwv+sLN9U2L9JcaVMlHeUETiXGajhVKcBJcgT6QYwlnGZy4FsrZD7m
ZeabhAboDbPRhG9IgSq6CY8si/6DB8cq6LVOGisRSd0M74xcWn5p0YG4XLUsYWbfsrw6IkFgw9du
F9kzj3wfL0y5BxhkOVqMivftBnUtmZerrYbJc/XClGsGSN52Xkwd6gZohBT8rK/eAfkNFNqTeUax
WJUG7GUeMa1EV0Bk28tOLVgR2nhRmYpM58K96XSPugMsayrO72jWAaVYZj5RisQEaBH1tSDJElB+
+ExxgG946G8lIC465DArGal/AW+lSZbf7RdICUlaNlBDYklUdQTxqfSURymZPlQ7sPh5MF5xwTi8
iF+dQKvilixrvHe1GwPiOayba/gH0TM3wlvw44hOhyVoQlrX/xK0lDsDXfh6BBP9112EYQp/R6pw
+W5hnwZBbITelQNbasECvsAh9ZdsHW6wixeWAb5EZiw0xVUQF6P7fbVePwXzx0aKh2hhO5I2aWvY
0GiZOcsvRIh2SAqA8L3gcwSgaj8bzQnbkN5TZSuGeKCE5Z6gNrS8iDCZBWCQJlQzkA4C/sa74WSC
W09/Kb5Iv2ZwO/Iebms5GrycDgVns7B7YjC2atBw4dQdhzamsACXTetUcrxJxkFbpZS31mCo2Fgn
sJQnhGtSjqzVrQdLmpo+5DWHtZMID1+4o64ZRXDcKcGKPrmGNCkrmljQBu+QVJw26KBD3wixNIWq
J5AH6OKLK8KzBvWhnsuk+Gu/fsBMG9zd5cSZqd5LuUycf9oiDJ4oCGnByV3ph8cwCtX13JybCLkR
XQXog+KIry2VhUcTeBYvbUtGhkR+9xe++cK9zzDaGtk1JvA1mDvpCz1+iHeHBhvYscOUuEXmRJvx
BjuNXBPaLMezZ6s730G5exIrKZYMOMAikMCBevlbsw//J6cdbezI4UaOrPpojpOaRe7CEq+sMBdc
Ti3eytyU5PCwsNxidlm1Sn1GHLJ1y3uHN+6DhQVPHEe/kv449oW/2goDCoJ2gGnZrZtgKn+Qa6fF
4e55XKW5B5L4VBt6MeYfdYEd2b21EEsISVlbdOuB7v+zBSsnhLN+UHfcB0TTgqSdGbjLNVkfDdGT
97Gl9fI/KEZYFWzAjNyT65f9xf4SouCmRHFidHPnRtFClGVgSpB7OmfvU1Eroc3gllUy8O0XiXvu
1qLipzGCMPsGsvTPqI10BflVz8xXt7HpGE518q11zKv4Mvm1VxBko7Y9dnzak/tguxijy6+NFT4a
YnkligefzVYqwcH09k9vxu6Ws/OGE9yuXL9TgGuw+2dOkGo6KH93o1u+vg9Ulqdeuq69QIqq9/cE
SzBUFPtP3pSggNipANDGVm/fjsMIbfuQwDLNVfwGAtZ4my/94pOAU/EsWv/G5x+ytPwOTAiCDFVY
Ow6NDA8sFbKpI78krcVWrSvveQOy+7HvA9ReILG5xQzApzLlvG/NHebG0JPwhh9cZJQmy4NmbyQr
10uZHwL9HOiUGuleukLg0T6uJJhF7CE2YtwGmnljGr4xlvVm/WXxY+0R3eh+x/k7DH/69sreGtpd
rrwie99kppevGCbEJrrExC05zZI8TVOw4t8dp3W0XGJVL/1StpxedgHZFpX+95Trbi5QgJcqPZbc
G0mhSPR/Tj09VXbrStTCR68mIWAKPDpVmyu2mw/+BYy4AmKVQYCwYGlXzTs2sB7XY0zApI4dWEtB
1h8YjNYeQwOJz0rPLekuCA+DFFAM/nyro6W4933TuXmceYL/4x4T/bzucA9PCV7xiuwcs100bArX
CYmKw4zn0Y3V6fK8h8USbrW1z+VAEhnH4YmFX04xakQUNx2fadKpy65psNepBE5vl2r+1GCJv61k
FD+MPmvM7K3OH7lL3aY4drJJJHaf64rcLFX0LR94wt4VpTSIiR/gsNkXboRmpgwKWaGmEBpvsKWK
RRKmA7XtqYpAI7KgV6PbL+DMKcAaw0NViVh+ACtKXKXNYnxz31BHqi1is8P5gqECo+l9YjeXPF8b
okNW3VRknqG/UdbVlBKlqV1/HbzXKQATU4AzI4idqDVqKk/ixxqw82MIcB39OPNLh+5Ee5Y5ZUy2
5BIqZ+/d2QRndUrBv2ILBFHXNEChgDu7h4+K3eQLaqyysTZaT4Ap1Wmw6EuZsBi1b/9Jim3gVD1m
dz9cVqS1XP/cpyfCOeGev5UhuxXbQYm0RSV8xukX89wb8GZ0R63g5oBKwWPYohdxvsza9pzzTo/E
w8I5wrruRldTpdsZpJzPCgwU7NXscVPRE3vR1i57V68j1FoLQFbCyGZx7n5w0o19zE5hRNs6ul+7
uIsose5iPBMhNc3KtyGOzDsrAfsnFqYx9mhMOoAa8jY0kVDZrwycjpCwSOqIE5zZLBkjtYh9EXlu
xuzEoNGZ0MOL3F6Iq2+j5bb9+/WohCYyYH5vi4lQXkCAt5N+Esu92ycU2LQbJAtf3tA9jpWYGyQa
ln9n0Hvdal7+R4+lVyTDGdSx9NgKLGkph1hSJiHddPwvLm8g6l5UzUC7Qm0ijbMMxWBdA2szz90H
BcEWyrffI/1UmASTRQGY6D1Op5qnb3I5k5vUqD0V1lQ+XFOy9eTVDyDDNNzVkq+/qvsn4DJVNdnc
8wqXIMrsgXKUOqwD7k1opx6xuY33F/954CnA5JDSqDgMJKgNpCgDA1uFkukQyXIbgd/teHVzFe4Z
hxMvS/nhR8BzUecsPTIyCV2m+KKmmEgnjprL929qmCLR+jEfOe5dYMYqKcm8/ziW/T3L4l80v5hp
ZwYQzUctvnCJyx/IeCJ87xNmF1d13iqZS4Tu+1KC5ZctIshOwFIkIyk4hJYobVwdy2oepKuINmaF
zvk10jXqdwIkgvC79De/Ns6F9SOadqDU4iTfhsbZKowxDtGJAiaIM/+6/X6zUtO3KVIE7DK2CXjk
Unm6yIPW0NZQ1ghQbb2aP2db0xsQoiCcHO6uTDvi4UqNvEJC7Nl/BWp9x/VCPMsEotCsYxgDG3yu
78dybDqzGxYGToATRElCMqYS/WDXlMNnMPq2Kzw4vDTosNDtUiHDup+kZEzKtCx4tPtMwGsFtHji
te8C9t1lzDfEowA6XZBe5opBdnqOeWJTBjlWL7wuuivMwgSC5CLLD2mt/2DlvR/wok9akwXXgZ3/
BLAD/exBMKqcv83G2dMN1jl2mN6Rinh2fAPRgaJx1p0EW9N8C9gO3/ai6IJ+PIEbxYhW8kok6I/K
OeR1c6NqRFJDOCHTKEkGWjEd61A+cSVqlweKSYQvhn8zEULHYZy5KUEUAFvOBkmr/MQ8eJ6xf5TJ
jDE/rFBHYVKuTbEIRb7bmQMLkqN6Qdqkqe8Q9HVgYHNS3MvUx5V4WanHDBOeOPYUwGc8E6VoQigy
/vCAb08Tx5EcURDm8xjtw+vT7czqzUkqqDuaMXuZtS34U+zgOSRp0NSKHH9Dq1JyTbIHtfmDLC62
X3u5Tm6/imtGoEtknFfz8LDOeg6jzaSpKqNgsYmL/FGuWawAsw5WAZ3YyNxYeZZnMbCYKW/2PLbF
Qh3nBX6U2iPfnEaMGMusfHJXMvMqBHKtPSh9Llw51/53l1X3Ped1e7WGz+0TiMe8RLqnMQBPUry+
8NBkEf1OTkY5eIc+pZuethzySLmqHUNek0ixNDtlDMPx8ieflcfUUpMDbA84h6Kl5OvVfTUJJ+K1
9rutx2gbrQkSqv9NPyhyqEXLGaLiO/4r4QBwUirX6PVMi5OB/qWwSVkwvIdJYuukn+Z7kuumYIn0
033AenavDduUQMXK1StflofDDW+/tQdbKeQ8C5RAL92D7pBJlGecr5nkNYQ6l1Jd/kBw633xF6JD
gx2nuDr7I5f8afsgnJAluUKuy8fAKJNCd9jEE9KdqhMgekmheyLqP3vvQguWMTKOuADzamp8wyVg
FubE1/+pZGBOmh7IpE+IJBeqBxOKDA5UGuKr0wMz441d5D9eM3nYJGFvENDZDjySCYzoIiTW++bp
fiHmYCZzdtgEW/pI4xGyCmPn6ySHZ09CYbHa5Eik+rtDff8eN0X1LeJlMsE02zMTQAkG4c8c7RaB
/PCoaAANW1b3gh4WzvffQooqeSPqmkDZlT9ggDoJET6j3mqCzLb7Xq193yNz5NZXbokLv9zrMIcN
dZ3HiPPoNIcLC7kE7LQzBwrvwjHfQx+sWi0dWiG2ebnVXD7S7BjPYcGL89z0mJ6oKnDAyIsxMUHq
yD5U9oDK4aEay7PNBK3dP85Lez4LvxSJirRHCxGJmqpcnrWgxoMFOpdOKmv7kgwfYlrfOqgGoMEE
897yhIcdhtc6FxJsPHvbRlBseM820n/soppK8j1SyHn9zsP9nnnUiNDtHd+vr9GFBjbNxu4mgBwn
dlhSdJ7NkHmkO91G/zOzACQmGGg6yQHsAHh3iGbseXgW3B8+fBK6IgZsNgOOlEmqslmL+5WuKvou
P/e5RtcCkGmV3mwWadOIVh0w9zuBQDou7BXbq494nks9gJ5JWglD/3HgOkWW+RY6ew5KFLpBeTnZ
FAKngjnI+yS6Kz994aJbRFPhpqUVTdr2mHZkGpbPlkPV8XekUq/COOzNQxGT2qCoDHImjfj+R+5Z
otKmhTtg2U8O3Mm1jrK1Cf3zthA79nWPXgN06gtT9Dd9J7Z5ALzgRbGOvg0QpY8Klw8WbwY8Vj57
LyrhMlnEd40TrtZgAvNwiYCrmC3rkxz0/E8eSn3xMcw7pxPOQHA/E7ZDoR2d+9h4xKdIyBlY8N/y
Qx+TCZyXqs7BSP7aN+At7MLsVJ06Mgi6k8ObELEquJ01EeAW1HNFp2yziKDBcdJ0oY2KpjAmYMr0
2h2EyP2Y0onVUNK7Y+jgekYBtCy34CRRbv33L8Z3EaXLmRa/oNNzlYTbzUxqMpi7rKqFcRCLwkHb
Iv0le5zMpJdy4VEbrd45Ny25lcjgxPy29JVnGHmdtcoh99hTEKhm9dtLJagqLlNd61j+NtSUyEpX
l9qv4bXqaKeZ8989UNgNOwO9QTE+h5ZYBr+c8NkEGCpGp55BeemL0PxmA28+x5i+oAUKMeOfMDa1
D1uHe6KZ03yLYRdobdqSU+y0VjeI1EHQhP9PouQm7gyaJpZiZ1M8cCsIH0HdnVf/VEfGJLm0hL35
zn+x5EYal6LUz0IVaOt8aXnAj74ZO0ViPM7pIsZbTH94UKHfA0Rw5ZMhvWVsmxZPBjRtmZkMj/ur
0MGD6tE8eGCavWFbxhF8JJlLB0P1XDTgbLUGmo8Vq4cbBqybMew5ac7Z4brfwF7jjehZ2zMk8lum
hFnFuSRIlQVRqkqOa9xlEbCHXIiMesF4StseB5DelkGeAmpYSIhF4dAwhCO5542l6tL+d6YN+5qT
rKlhLqzhqSFKWvzaBU5i7VXXZSm8BQclUg0kWNPI8787g0k+IRrG9P/VLpEsLSYD+eXF3jGRaSYM
IAeHGw2ZflTmmuhLWtu76/wFsQ7gjtxhtb2A3hAXItkdOjA06U082PYW174R27BqL93zl5LcJIb/
TuQBT2UJ+723WZoOPvCcCEUxPwbStzGIcD1Y+xKVnJTGkwghOPs4a/TyRI3RKZlv+kQOOgZLrW9j
56NOMwvGO4emS75D+rWc8HG1luYwi6SSKy4lF6QzVCRG8CVgevjtEP7R+MSw1z/mKi/N6CZhSQeo
NHInJP1X/muFbkgYhRA1r8LCZi+9OhRVxFE8xBWweri1+hBzflWVIGoVzD0nKtlcC8WCxzktzNNe
lEwfdB6E3nmF75vffs/jbZRTtTMTUKw+tRHc1nPKAAicrh7bqjiLMjdLPR9LNT8w1Vwfkxe8dfTK
gCTqiCC9uQBtBUZvlCrP9rmGCpDl6wAWxN3OpyVesRfhKBUlyGruoTWkaA7Z8+sNyhsDZCHfGMG7
3O+YXFUPw3ku3EvOjf5EL6JFaz5yVrjZJkilFntppv90jm3kPDOEcpjfbvqwLJy5L5EkB1KNXvk8
5mbXm0VGGpXMh1tpTHt4cXPDxkUK2tx/i6pFqymAqvxwYgKlVX+hjaBL1LyKCe9ERDQCi496Vu0y
YRsjFElXgmwoBbEAOCWwX0zJcfQlkEQ4fCtZVI5XNyLOxkOPjnizV0FuwzrnDBUvt5VOrdbS6GOU
t4e2YQ2vaiaMAzx5qLWMREsDBUktfhEeN8aP+ma8QHZBw04Qz2U0cOiLaLzSTWeUH4Bsug8WFJQq
02/gS4q2dALwb+VeEhlweenUjOveuJjgjF8kob4me83CBMHVmhHNZahXh4dJXtk6o1IdKBA/qrxj
jqgXFLZQQa9ihkFxvzYq97GUSBWY/+Eka2MxjppGfAghoGupWU104NrVHSCClCcxLuns5CGUditG
0cmryrL1UFZz2IxoZgml3cE9D5GrsfsXJLG4/DuvQ64KZUziKyGhisblDmFz3GyqfLC985VUoNjH
3c6xce1zTgb8KSQtzsmP7LmUou4kIkwMfDVYwDmY0QLX8oTs+S18BefWCUBWZy/07wsu0EfEPmMK
IZcLPmVc1TMZhpM+dqoPcoROFLPQaf2AV+nHVAp4I1tT5Yn2Mqn0nNXk2sHhItZqYIRxg2ouW9VE
u4D0plcQ8Njrpoey9Np5UvY4YMprhLhR9sf5sHs+JwYJMHj4ui1VE2FJSV3EOuhKzBOi6A8sUhjY
Dxi+nhiNMM4iWQpKIkSS63/UjD5Br3TeDoTX1rGmoHy4zpqlMTmgqn+iIp6auawsh7OxlrU3l7nQ
b3XDDedFHQQb+kc5uJeDDaI+xOuBMyLf8lvtnpbo8AtN2eyfimIbbq/sMEBh3VyHOtPU1MfKVByU
09N11pp5BQeZClVr2LQaGn2XT/sQC9fJLPVFyGkK3Y92Gfg/LH/JvmOhmmD+Lf/Wnu6gDWhFpHMT
wb1SKjVtki2NrBsFCpbtLGTigJU/ymH5Oo8n7IXINda8SBZS1IzQ2jgwd/Tpk7VH6Ut7rr6msNzR
MY44+C4Z30jFvYM0VFy7tb0iicpL/mT7cBk+2mkAhxUUTydZbJmSj9Hu6PgemQgi3p4/u4VZlbJn
CwkGgO6CrLH04uCfHilqUgAayqWlfMKJRzMn2C3foAaZyT7NPMPbIrXD0HRMal3yAHb3CWpPJq1e
6ix5hkIdcrtcDCZaVfUeAjF/QewHWqwgIn/OBC6jZ+19kDHBjnOXkQU14JJxSInDPCpmWnl0ghPP
pJXrHfcdmJZLYq7xtzzcTowv3Sx5xJvxVh41pWIi6t1yM8tOigqB/BR+/0QgPi+M5HZtQT7UqgOd
hkkPOgUmfuNQqEDLyO+reWS9D4jVikWMvGYV/BdjDYP/zuhWajSwZ2BAnA0bSFqwLqBLA5Czca7P
TaaxNO/4A7u/r14fEgElU7BJruVg6OYR/zt+P7b8GSQXu2mb/ByaIsI6hgenC+07UabOApG1bWXP
IE34moC2k+M3xAqK+UphAJ3o4KrJ5cgyrvj96jpeCJCeDCsFdMfqyP7gLPlsMhebnCvk+0WF5eOc
7I2g3AKtqj7fr/7KBgUJ7jNwTr25QEPj91yijMjfk5J/hJHI2XUW9bJHJWNuztLhT/ohwHHWWpB/
3FIyY2HlZF/5WtH05wy5tzU2m3EjJXNxM7SQYZcQ7cBuaevG+YMbz+uPMnj84CsGImDH6YnB5YhU
MSKPLHBKO7A+XOfgyzB187Abub6IgqCBUYv8wP3qmRaDynVl5DV9xOF4poI2aXRosDuKpoF1Skgi
oCUPl7PSZkeYWpp9GHQ6eVzbpgNiKdpNBJSVuV53pnh+7kQFqFcmyb8drVDK5cJLKN1kcf5MdKfC
idPFcyo8g6E77BfLqtvBw60EMDLH1YmtyB+Hrt1+m5GMlYFMFs4UDCXFWxUJUm6HhJEcIaRpraOt
zoxeZLgnDNoMcA2WcUvWSVZvz6awkEtJ7TfDJu9CZHofZHShUSQIhp9u1Qhlgc8fdiVFD9ezuG6e
Z+6aaHkJwVTuOhMSWCo7CZDkFw9IpLAsKUelB4txvJ+pnEEppeStqgcfN3VyIQtXVC5gzio5Bf+z
ZC7JNkZmIGrMaZjbulAaSbZRQIGN83EkB3LvPB3CD0isb5+3Xu2iNsDNqkdw4qoJnZGIYt3nHJ0S
xTlbIVVtGhnnrlJ/UInCjEarSC5ZfCEHEgYXwQ0wBbAK2PlhItiWnAPUjMSq+C4A9uYaYn6nVWic
srSCYVZpM9yCCbtSLD3qTB7JSHI+hSDLsTgrr8qyGJP5y/nMfP6Ztgi+HrykdubLbIKGJIEYU3+N
rfNyo2vUrj9igMtukbckXn4R8vKVYIiWCZXHzV2KopbiDos4E18ncfFOCdBoxRpSkALSEv5JGglA
MFv1QufK5jzDmj1d4tm3tnyJBxPw5vN5r7ab6OOFb/F3xFzO+nMyI3AkbYnji3X8tuSKMWTQY7iu
43k+ynvoQfxre67ODNpBocoaSae4GX1334uvJbqsJAHSz8+I5VYQUWt95pOIoaCm6+XMI+oPsbhO
onk1qobRaYF7GdwJ3C055Zw3qbixQQGYVHsD2ohtxLYvEpJ/XxZGfu5Zq+4qViPS0VYEoN4zJ1gg
l2ZugBuLyC5yyy0uxFAvZWgUQoGpCQz3IZpE1XZ32ByQYrKd/dNN5fQF1V0lkZnMqYxmigxu+VpG
NFULWQXH2wY+/0c6ZyRSde5O8beV70A7DJcPzXJR//VZJA7dotCuDJmNw6lXZItAH3ns2/Y/1kio
yaIZHnx+h9xGCZ0m+FN48aa+9UexJXYgmOP0RWBj2ZkQaYO/nJWd6FJiFVrEwVMqRVtYrQX0YbH9
tGVL5UENsJZKmwooTSBB1Tc29fzxTEGxWH6eJ1Q+oRCiFXfS0QXZhtAyB58ebxck5DMm/3F8Ozsa
+gt7IEzHmj8fGwVVKp1Bz1FCqlb22vWRpoDlRKAN7u3v3fGatPBvtnP3CZHaQinB9AFfALXafd3O
CqX+d+l7DCqS+UnzAOx5U+XfogBWejjW7tr01uGj8NviHodFwyCghC0P9RdbYXL/6mK0VESWHOhs
HXWfEcG+d8dntVGoMvKV+Nzk0VtuwEBUNqwvYLeuULZXDGv5O0p8uVRxO4KpDXsaFvOPeXnMZM25
rwUUSsGaPd5lhuJvDcZCdEruyM9S/p8uPWSHhzE6XEuo5HFCQgSMK8r1EaeDlxP681A/vpuQ6MM0
7gAlsnUiDNrmAPOXpTauo1y5bMeoU1vcSHpqFmbeAIKJW080HA6h/at2c8js1V0oQ6mLElJ1crHK
L/TAu7QlWNPy8qYEOOI5u+O1mYrvONVj/Tw6Hf7bi3WptTDn3VimwrB6CfRvIEQPuw6j8f96GUWK
jYZfJwnfMsjp5yV/1Dmsvw7S2uep8x0ZNzqzXcLPjLD9ACB69o78yPxxKRlcv4r8InlPVKtqfN0v
MFuA4QbA9hMTCiWwaY73Lic5wkEGYSvVyunD2DTxa9ZC6V1ya+Tb1By1gYnXKnPu9MRIq1EfuGqC
WyHMmft5g4UTXBycGSpuoJe6i8j4eXX6LskmTQFeUlHwIVv191xtioT9XXGaJ+/UbSufM+l+CXtg
MZqes9yxX62eQ/QOCEAiU0UScp8fZ32fUAulzuKklE8hmc7iU3yUzsvsVCyFigA1ATBCU01JDQVG
cuGC4g7Z9Npsei7didGWjHk4IaTSz8efCRHUc4tghmwS0RK0hzF7Xudj5Py1q8jAXMjAbOo73Ncz
jJl94Q+0MtuAiXN/iqEs6Y+glJT6tCFsCNmrD9l1Zv9MW6wsLXjxRQUwCfEVDItQ4T6q2cSIaxNj
noaGWe+GZnA8jiYJxNiz8ttMm1I3CKyaR0zQx7mgZrD+UTEIR9WLRMc81OktjMwKejtuxU7icgZ+
I8U3tuZHi0IP6t3KoTck3lEi5+a5XjEErQQCsLQX12EYVkL0e6nUaWnPNUDsQM7FOSeIbuXmZGQ/
8frMEig4nXqaTS4uvZRkofTlcD/5vUsjE9nC3640hXkCZuFVAReIVvddsOlaQtFLjoEmDYhWSHhU
X6/DZQs5+YGMhCd/6ReueXvLJlWrmIj8Gn4imH1I2RFkuax6JrbVzKi1iF1fYUuhFh3oH1HNCgOv
5LhgxgqfWnkOGk+WyPfjHPaUiHS4bRgOk/YF1rQaqgZfkN/EtYCg7vAAFZMk17GRhK1hPHboZcDN
XW3+6he193bw5qXwUISqlAOahbO2SC0UlReHCEJ+iD7zG9nnFAcQF7aKJAG4q8q6fW5qCawa8sZ9
IVUDwrP1mRDnt0dNLnr/LkW2v6NgoA8zOEC4Pomehn9nGweADC29fUnetBgQci1caYBbqhusIUSE
3aMDsbXxcqe/y1rhwNmGLy6qzFrioUVDIFIk8I5MNlIzSNBm+elUdL+EV4dIjh3KKq7cf8mGbpL6
SmSyoCp+u6/jNcOsuSqIKAsyME6KJsWS7k0RtLp8SQ1uRXBonIwSGbe0xJQCHahaFZaf35bXRDep
/XLlzQ2+jsRiYC8cB0PwswDUa5P6ISZM02EDqDirHGst/t2LVU+2aIpsK40xwqfecTRU/CqiYSyh
ecTVwpSUMexa2QErcl+/RxB9z+QOEKFAUswSBPtvrA3FIaKx54nAIE8vBnl1WigiJoVT6jldYGn4
mzHAFqEAU3opJlTNxYwz6uXZdUKKlH302dgA3H20TKjRxskY6cVggYMDeu4iTTQgaVjK++epl3OD
gzLVjfCadybfFiGLHsGO5KE75ERglC8Yxy9LzdmeSSU14btpiMHh9BUmw9bwiam/W/AKxQ23ww8U
shHIyaBHatYbdtaZfJ+Og3XFLkkNH3od3Ayk6WLiNjoThUtHoV4JA8jkd+1g7kMtQw/YVOy2vxLY
Hhzy5M32HeP6t1Zx+KuKGi+5067aUPYplAf0x+mRcNIfs7dp9F0QoytU3kqiU8hh3HA7MvWmREI1
4EyBBUiUMG/JTpTlZqwrf5v2/76NKt8lR11Rrp6K36vlMZyOmZJbTallhg++kvYciQh4TFc+oORI
nWh4qknZo45Gu+brB7qxyILjRjYfhMyFkdgzLzwMPdhBl9JXoJ2I0zntkR8Kn4yijMXy4Pr1ekDu
d/+3cWLYa9DB4sSVwwpYQPRzGq5fXYuFC5stTHh4VvRLlIr0XkD3jWzV4yD96JDuGglMWgXA5KIr
kb+nbd78RoJRbbuQRNK0Yx9+vm0iYJgPE2vwBp/c5ftOtsKfb2kBOeq2xwn9TMXZEDb8SLd5+/e0
r5sP0LFTF+zEfhnMDrjBW1BafHnBK0G81ZyNvNmmxrW1Ue2+RZCibiFF2zufKgoB56K+JaXZlF5f
NL7FMu2pc1qX1DHOgy4TcOD6b+U7fs6ggM57m3z/XqQGufvOjcQ9bjI2sPx7FudIuoWhDSLCT/5f
XWT593bHB6z+/dtW3HCfzpfMQvHIuTkIUlusJxgLP3Lne3cqz/jNjeT8T95/FFdinp+m41zGi7ma
F3kPRjOJRgLKhzZONbXgqFT63Kv/gVeRkbMfgXk2GPZQ4ivSaa8zkBaSb0sUuDg660HXAyTZ9yN9
QN9hVlDHomBNpOTzeiYblijr0U0RsQPQRnjhWwfw1bXJhjM0GRRwKwnjJtgmhumT4AbVAipkcR00
5JzdCURA19ayF+s9FvK1cqIkW5tW1geX3n1/GhKBZHfX9TefZwS5n+xBA/SrBKe0WPuCp0melWZD
qp5HTdxurx2s8KiwfwnToTJ7Je2yVZLedrUQ1/5NTTQIpZmd/8UG83RxSYiJ27gC7oPeThevBSP9
29Ev7rNTZu50rfJ0fhvyzIiaAGAVymp52q7+9As4X20UtNAT2kFZIzgzrtVAFovzTI/OLKUnjJs6
HQ0IrRYZ4wOLwRze9BWxMEsizIfGWjTL4imy7WlPuxxSf34WpsSKn3i3Hs4sfVpxZ5ENsUyxcnhr
Y2B8iqNAoybjHnfVCo3ABs2I0JKwk6N4NwdiXiECsEjGgW2WsRUpVBLUiyN9KQdR0qp/i1LAacmP
x0MxQ01Mrapi2DPeva1uy3My3wqJjbTHfwdA++Fh8rbfszcuRVUZpziRr839/VAPMQaPcnuUVI3w
wbDJakwRfBdQcSWQrzh4opPxXhJMkmxqBZEc4wJxLwUdkZ4dfadav4Hu8/g2iW4U6uA4zFHUIfPb
7UWn+Gs2uzne1hqa4beJCyWbm4Uf3mY/5IHjIcoFtuvZmfTB1DaGTyEQAyOroHjYDPrNre/csqk8
+osZ69MJryVDHBZXnaN5TmtQ/M3WXSQVZDJSbCVSmwXP9cnkHruELSRexgPuNtUSjndP7uAWWbiu
x0ZW/TKE4FsCI5s7mDZ+DFEgSkFaba/pmephWuxMWp/DArb6iVtY9Y3NIUmxnsjRXk6hkmiE8TPH
qhSypgzY4ZxSZwD6Y+CGlW9gRAAU45sHhEV350HwOCzTbyJ59cBxfG4yystu7SKZofv/p2zpYfiz
BcTUpl6ZqFZEBhGvH+GFbet1VGceB2haPkc1zO8QQzmBl6vfSCXysx+4syEwycDTNvBi5N2bvTAq
u1Av9QSZXboLWkpO92iWuxJFsXZvNId0vjx7Z35qzAePXG8YKYHYd86Y9002YCUDPl8jg6lA+LrZ
Kln1qozYhZhTU+NAVYC9NZB/gqwPWpigSM+Ag+L2aJh4WBByGRmKJK1KVqlHQ6WThOEVl/3Q+6oa
151DGZ9zuKc+2kajeAjPeCyF0FBEZqdVGVd5TqIFUv/N5nubqDqPAOpiQt+jy224FbL7xgsMesdO
o0fuH3Tz4rOTJluwY3nO26uzw+Cf3+HsBdIMa4LGGhWVZe21oIgDmzzua5125iyGc/dB+x1W7mpm
YkFMHt88z+X1Cl0O56lwuX2YXCPefxT+zjO8x1FsV886V3Jx+kkkWkEou5/A7QJr/muJ+4/t62oI
u84YPaIceQIgIsWk+pgMIm0xmsCkSHABAwDY5pp2hM4jxwhW1tEoX6iyy/XRH/JPJ9KoxTG/iwiR
PebNZktkwRc4Cgmqj5UeGUpVO73/vj+v4B9xi/VaqkdVpUXWNiSeSzKz8d1UxcMwiQgy9NZQgoGh
0LNt2avFYNZhwayXJwInzk9rwwoPyowgqZOLXI/j4Ciw+p7suMZevmfHOhuRcqTTbLYYANorY0K3
7QO76spSgXyWDpMB5VbqVruBug0Vr8Bwa8w+XD/inPn6B4VW6aX/zMIUJ8p6QCuADiDv88MUYYw9
OLB6P7//njhw6pfKf75N2qQhDpebrLr1tjXkT4XdA8pETr0Oz0fd4qDbOOi/Bx4C2Ulr99X8zPys
jpLxfS/w3HS+ccbeMJHz1d1n1WFBdOor8C8OHRepe+MeyvwRqSa5ZrMRoMZUDvPHoAJiRT24/c4+
9a0kNa1J9i8qR4IAzNkPYypIbLUel5ZV4sktcmrXFNOC6Ne7Y9bRW5ZMvqMa4c8N0SdWKRgbqeKB
3C4bFkHu6kE+R2Q7RtmLy3PpyApcYiHEWcFA0ZPvXsFIlztYHXC2SxcLLNS354LOXWGXLMdpF7he
JATVmLMhnV/YqAIb+njofP0sYn7JU4gzdf9EJ0p6/l0vPDZ1OjZpMcPdkW8XBhdFIpUt+jvUMwBW
jgdjOp9bQJczKLvndjyvrNfkv+BRP1GKJ+mn/HI3RzMHZUhCCai0nY9jdoeJJMryR5S1Y21MhZj/
lDfFnGzHJpg1/QVhg8PQ5Sz8SZR3uDdPgU0+GN1esNuBtc36vKHk8wZMFATm1BY2ciM9O+igfmvQ
GKRl+ITtiSJXyjAzv2jyleeXAaLbQji6fVPWFgfCN+B+wfkymfc4CaqYYpZ98ENvvbwzOATOT6uD
d7VAP9y3qB5Y//e2GeEhPju0/dCu6sSNYktkeRTfTdU86KEMn3ACUY9Pi6kja+HAusXE5UVfJhKK
mtc0qLIjMQRAz4t+WPRWoI4seRsV7mxY/fXhRPUew3hYrygrWx1DNNgQH4QS5CiU55qqTqHB9hCc
Ond8P0DdCmERqduN2tVkqYs+gXWZEvTqhyIlUwGCvRdwh9F0cu2sd4Lo1XUsniWhP80ivlQWcTvx
FC7Ha3PBBSuYvSF8MRlPb5hRzqD/ibT/Pw4msZw2KtYv1UWpmSgZpRy7EkZ8E5c+tP5gLM5o/EM3
b+8fuXwsZSJM+mvDDzJRWJhGuIvcDKa6sHapowSWuHK7ot3BpUT1vzztKRd8HgapIbDg9fKVFUP7
PFrTt/BdLjH5knGZvYoHKTQ+4mOK2kNXn17p61eDohYTRLJH5ItI/sGLP/hdOqxlsoiBZX8+wVNe
HgZ4zvSHowvWnSz458KFGwA7b9IiJ/vPjqQoK/87LNJjd6qo4r07mXKqw4pCUdPpooHGiIkdm5p0
LizrWazsHpv0i6Z7H9d9N5GZufvYjgdV8DriOkmLEre/9jIiHdW7WP4nlUJ0JIq74XR7tso+JE7w
+f8b6sVLPXikeV2hnNKM1XizbxbPE5GxhRhPySqMaGCsoUi4z35kPq7Iglqggewj5nG0+nY9aGJN
FNKURkQrNZx67wNyFdtnQcpiiZYUvwMaB53zE2v8w33QkwD/BGbbyPkfHq7EH6DclaVGPCxIIjx9
OzVp8COVTzQr3D+Hh7cbE56YhHbnKkRtF6QodZ+Xmhv4HtQ6zFxwrztJNALbhF378YuMdgUpplPq
2zSq2rCewdocGTSaZvAIjHORgNRWN8P2ukBmIW+CiqUye0dt0CCnNnx2m8I87+3ppypaodvrXGg6
35BGzvEFs0AOjHV2MGei4tgOqamDErW3A2dijcBaIN9+iG0Ibh10v2y4UWdM2f8Y2TW+scVn/vHW
pmLlpvGA3bPdIphjSTUuaah4iVVcIqtxAgVYZxF+1ZshLU/6NQsJ3cHtzqKZ2uJCNznj2N7UaLfl
2Flw9MxHKhLb9/9Z0Ic/vjrBueAAc2MX/6mzcuftMe6P7UYrnh74w9nm+DCZ5ps+n4jKBtI7Pg8+
p/cgTEFOPip4mQDv/zvrfY0Yphg4rAM41qEYbeAx6Ra4vFQVV9bcBlrGd6IeQp8hX4pHJtwSyuTL
FtHjbDOZqYNVg0Vn1/nolrfsvoSldugkjmCZsq2OB7q5mKMkyzqq+t87ylu+cvSUy/JLATEwGaMr
FiWQDs4Q72ck/SkEjfVY/xAkw7p2ORJGwftGUdKpU6PjGmAXf8OuOZ8OHLoyb/exTvC58Vml+6+R
dmBTdMMIuKv1WJGI9GkeA4Tm3MjBTH4YDBKLP+p6K5CsqmemPKxL/6jklDoxo1eV2BR2hEKz9bmz
Ib6XqNg2RsVlxg7EC7skuPkUyicJah2jLXOp34isdOcCD2slA/1Hdigx2VD/wJqbC3t944RWTY0C
Qy1r5weKmUU0+KMNJQAaR9etcq7tipc8QGZRuQhewzArjtvcpTMOqilk4qcxUeYm8OHOKjCtGroD
nzmbda4/c5GP8LdI7qaJX36KmskBSwwgSxJTZWIAkK6H+C3h0wFOLGOX4/n38a2JN/HWqVJ39NI3
5H+JJlflUaJwAgdqGiqlHULXKkExV4gWTwhW+6Ubx0Z7SNwusDgtipiZzkTytmxVk6ImUVWN9/4U
UI06BymTLgnXP26bg1wLtqT1lhrxmWesTVfWT+4DukhppcT7EsLys3VfGXia2fLOoSNIDwsM/cQk
QiBhdSElhDdhMwEMpho0s2k6uoBY1ZexnQTkE/F9W6c2/c/OOvlZORqXvg/QfBg9Zcjk+2TxDqEK
QTHovrB7sKHWrZTTaTJDusXhTBKleYf7vcNrEM63zXgiSsJvBczQcucdifOt6UAsSt0Ph7C9W7f8
IASfNADRmXhAr75HVNGmnlBHQdhtUk3i8pjzc3VThP2o6pBv7UmakLcblFtJDdzcyf8jdoxlTrM3
E71XJ3C7Q/kDFBUCS+2j/xyvZRjC+5JMZxLLE94p+PmR049dOcGLQdjf/2C7yzHiRM4pu8eaLb9l
kYV5HYVTYFBPzAmgF+ZrxdQHZ+ePIJSXP+2SqFNhpOWH79IPskLCnjtMHZfEKg7CnOfxhsgGYpx1
by6i9weOsH2arLNiKjFEejBjBmcxCfo0lDOeNh1uhPkRCqGbLPhUfcw/Xbv0xsTSlNrDpcV1NPjj
USin3G0iYIPnJMCz2JmPet5wk3QUibLlj+7dAq6kKaG0aigL9sUOk89DZr1s/33K7ujPcA1H+L21
14gGHBsn0KhAM5IWGgFvSo3csqg07STMCvzGOTE+bgi9T+kcsVWGWRqsVbE6OtyPl9acYsmZ9js1
Lrp/tOL5p+ujjBjZiYskWHXaGLg2wsnuIbJa3R3NBFBhvyJtyCr/eq1d8xyYPhPQeES7iEI37lx4
gGgjIwayD2KeOGARUAVRSPxBFpBN/7t96nS9j4fbZ7TNKWJIy/JuafRKVXiHNizyzIDlfAioKEjS
1rs6wu5vCIopF54pWFdOxXWOLsXJ4YkEKlhfcFE8dnAP862yIjNWIlc98IIQYWebt1MhpsrhGbRK
/of3DzoAPBTaRVUjGi+1diQ878JAlViwJ1xPEQss3cF8ghSrognIP3hO5+u0aZySWXpJuAn6NVRa
C68c2UgiXoyBafiB7SHxpMWDq9tTJeGHJgzb9LLb/EJ6Vyxvw40hG/p6X6Hntt53ll+JlvhNRw0O
BqRfRUmVb2WIdSOJ47Csy02RaJPphLKW5OVH54yhHeTE2eOkc+3NkbUHtJW5TqYz++ysx+D1T+VT
CN/B+MYWpGHhdzvpa3TIaoRcg3wNEU1sGGSCNdWNc6SF/epCbl/f+BIpAyUbwou3CgonfDWLzl2C
YjehqTH+FmsV6PI02lT4tSvTx0dmmYO5mQCGTeVhtTJGaGfK0kukth4rno3qhgnmZLUmmgS/6dK8
TOFZMxI6NL99bqZyKAgCUH6us4R4cxEz183Z5un8oQBOMiFOZeqF+60n8+5ejaDnQB+H0h/a0qmW
+Ql81OAeEHMJxCRHOleSsMNHL0eIoqEOkzFz9pB3U2joyRR2LbX2thfn4xDlrVVITQbe4+NiRbBH
plOfE1TiOlwPCKNHvMD2hzV4gbuuBIlyP58rctbD/qH8RLFRYxzYGSgURBlfWTT8w+VgD8LJ9bpH
TFAZNO8qQQ5BtNSIL+5I28EjnsHFDJsgWbUon0bYpgST3siOl/vkk7ewio9k2+knVUwkEO/Pl1ZY
QRZZTS4Tq6pDc+CJmbaV2MaQldEWB0ltgL0H0bRhSYlt2MxISoVoi+2Bb3FBLoiaIRFb+4uQlzl2
0V90sWdfsubfHb0NenW+diKsofgsBw2FQ3ZJb7h5xcbpA1K5MESUM11cn8rv0o+KKA+50y6VdvXn
uZLis2RXeGXDmdW2+VYuS/1KLk+irwxUJsgqtqHZtAAh0PV1J5AsCcsNR26jMLcgDrVEMGuR7pZT
e71ijp9VbuuRLfuVDWtTQcOH3BHunhWcVlu/VLaPTlgjCGlvZ5R7PBkKEDszaq8KRYewa4YMlhm4
EZj7iV7HhfxK5JeM/eY9corkYjsBrlV8y5pm7/CkPEksKT4nQx+3fj4tGw1O/tADKhJJKs1v/UZO
A2wOfrybXQ7KZ7OepbXrWWZH5Otw20bh2ANWg2F44Rv0zcp9qNPdxU1xLvHicvywMpEhJ2g3+ZpJ
fv/4WiFycbQa004mmz3MOuKobnjGBzFm6kmEhDJWrMPKsqGU4zyizCwnzuYXQjwhoGIp0JfrZczm
XTqDM4JuvDqstR+6kCjDT6o3s85ao9t63aZohUSbIi2BgfgudZ1DC+psm6+m1PsUEjfq2Vwk7wsv
HEQ5IZIIx5vcg+WBIz4yP7C6Qc3qiq4Kha7Va7bYBtX6ctoAn1apBHvSrQyheRYwUMwzewC3rzvc
u3foqOQ/mmS5S9/zhGocR+q6Q7CoHhrv7edFl6XqCFMohXQZH0y99Ah2e3V/iZMAobAE0VnbArar
XVQ3tIEwTVdXZw9Vdr5X73E82xsRDR8Anl9H9src+CDgaq32S0IeScZW2d69kVQtfZIxJ//MxI8A
27JENxMEHlRHD/nUuHGSiwj4p5E+m9minOnt+ymBWL66PN2JmaX/h+5qmtgwNQVYnWP3usaUehPB
J0PbrdoHnrsz69v6Gmxw0IrsOW7UZNK8Zl2cDAqq35xJt0blDx+3tJz0rVUGJbkbVKJ/hwiDC8PD
odfFd83zn3A5wbc/fbfdxlUFDCV2pfTCaQb+Xvl6561dWBiHr+lrzXvGY4iXWyd3T4+A4XO0QbCq
reJxCbmn1ey2Yb913fTtOhhgBJlTYAPPRzCZTlcmbzndCiCZP1xLP9WL622jG9rTiUG3R849W2bo
dsGyHOIUVu+qLe5sN0JgeQBfv+4LL4lz349E4VBGGnckICLyVGoQNcMjKtCyob1q7CLq+BwVkGJ8
1w96UhJyt4DIpSehi5UXLpWUHdHmYEPE45HGfhBxKf+BFFbpBjc+quYXTwu7MOZJfPtuPZ5igoCW
1/0QJD/KNjkxjrAJSm+COIcktp4Yqnf/lSznpG0b48ew+dqZ8zCQkBcPfgsA05V8QwM0rXHmJsFT
go2QGnHURGT0h7O3+39+9Gxgx1e/YPWaMDdjkRKkT2qYm/CObCwIjsAZkDTr11tGx5K3zt3OZOcu
jlVPYTNY8BNlgJ2iRBhpsImWBOFXAFlgSk76WDySSstrk3e56Q3WUCEm6alm15yuDSfPb6BGA9qo
mVMyypcD/h6wgYsgGlZnStnNkBkmd8NvuKNZO5xs2+Xbg8jl8nJDsiqBay2yhspQg7MztJUgnTwi
redVE+yt436lYieHA1UOisUxrQZztpMhoKKt7iZwSGDKUql2VpVZ9kFmrY1ORzFFQUyY/HNpVNdD
NkJzi40TQaLCsFUi9gl+tyzIurKjhxuNVr/PYptW7v5aWbjh4OESUDlxjsnySEGbOd5bE3l3USXk
SAVCqnkxFcaJ1XlK9IEoMfHWwWJlLmTuQdjcQzGkXau/DGvXCgv12paiww6PXKgCdI7ZBHNnH5Jg
MKzb1e/qbYBzTsrRKex+8Nc3pYDAdQY9StBT1pEyYvjPrA3IEc5t4b670KUrOp5e+ZaFaA4OvUUO
f4A1LrtSV8l2zOFWhLLtLPxKc2dLdG6Jka7SqzW4jiM0aRXhuuSjF6PvpLENPf/BNURVfO4K05lQ
eskdvvxnrlu5jDyQDHW/EXG6E7LALl2VPef6W7QR8I6iz47GQv7gCHqs8K3g4dEfhVYqd+Vipq3q
9NBmbZcu3pDULM710cid5usE/tvbyOYVYlEyNVp9ZIQYzndmRoGbKObpyAROGxSjG6rcBfmL+Sfl
8bi2CQibAYb/7R+xcs190RniwGmaUBd+u0ai3pXFL9jpFDgLrNhU79EPOZ70dLMdUnJNxOSXrY1Z
T3EjOSKQkbpl28P3cYcbq/nLmKzs8xym7+QSh0JOlPmpBUcu1Zk0fm9emJZGI99eHq7oN/lGF2Bi
NXf/vN5PYm1eyYVf4EMR1LIyGns/H45O9t7WX708P3mMdU13qxtvR2msX/TUh7D0IDfINLJWMykA
8FqQWZbvo+z4oVQfGppCFXZ6fzrBF3G4L1OYLeEP6EZhfBykv5pwj73aEdsyNZ1k5/SmMVWjQfBz
E7VcI1Rkzkz/jenZgwVtR0Bn1MTTsY1DrMxmNbq2r75797RnzgAoHgUVcXYmht2Akv73ZTn+M06B
YKg6VSrtcque6TsGmD8rugRWhXSOQbYun6lCJY3HwNWRpBUwdwwdeCoj2CfdbM5VvUI6vTW9D3C0
IWMFNj8/awFL9kcmTPlMeHog8XLPW8w7JRZdtmjt91WtXuK1Kop8CoFDQQS/E6kMGcoCDc0c9Ixs
hPEr/LnlHjQ8oFSE/MdHvkcKF+x7OM1KzkV3jbSnpidhfb/rtCrEOmW2ybHRBb+5uSZLJtAMm63L
SaU+766ThTLQN1NwIS78ugyXt3TfZcyLh52fulEtGZXIfY7TUYi1D+cha+Uo/gY402n8tf9xjeFk
RPIFDp+71VJOYvzR6RBebAPAdEfY9lR7bo1cPNfK95DPhkSjSC+AOff+SCbH8HcNFAuhEL7gXHBD
22/6EkAGcxJEt+Kcz+Xv0orE7kPx4y/wnYWaPHBKq77FqKF3ZyNWPNfeVJ8nss4taE6SaatPkPXA
dqP6Q5VkyIMSXjXJUCZ4AQMn/pg1PjYQY5ktVWZ018Dk7/zKq57KUTIMVrBq6cRrZCNSZV7n78nx
o3qTgswnzcT5hHr+iOrTYbvlBfWRI5UitYyj/RI7okspLRFyM3jz/QFVVIumRlrFMH158/G6q7hX
QNhrT1Elcokyjbk7Ry2+JZNXohjw9NnZaEyN64+NdxxYokgVovJhAPkNVaPO4jVCICHEv6Z++/NM
AqxRuKSCEVL2da4eeP6MLUfGEnat8QfXPvWviFbK+hVIzk/w8yaNA4k4ip6mS6sz0CqvBdwbL4rr
YlD6quAoMfM5xMWd8eChic4JQ20/qUhZO8K2MgHkkcvblZEUeReJRtsU67Zo5Bk2WHrnvIhViVH6
3Unr0bn1Bd9P7xHqeQoV0AghXDgOWASE9hdqbkad6kuYShWsfcn4nH2Ehu6n51dIERRAhJY3dcfg
JDTgE7DrfQ/C1lMSpmNqUnGrFyjeAJmGsvLt6w/mvd63BNCxu4h2IDTFdWwNyC5mrONTQqLjsRrR
MsxAN4RBybzbiinaKG8SNVQRDkFmcu2rUiQN4/hpw9qGN9E2etruM+vytAwv1dnQtpvBkg8rTuvB
kSYSpgzbgW8dhGsi6lgkRc0wDsz5oQDeXkQM8TbcZUQt4RnMRJ3AxH8w8iDF6CYMwbwCviGDyt0o
roRN2d4aAFNKhOjzNva2lXrcmBOWnxomq+wuofQNEKxtbUArMdDaeteNGSDyMNrIMKUp3m4e3QRB
6Gt7WkO1Wtmx5hXDETYBqCPAs8ZZw2VhBfBJc0N+TpS6BF3A9LgTWEdMFT08k8LVEJA84C35BVCA
dbnww01f95MBHbhKIsIQRr1UdzQ+Mu6egsOBjy6Wzm8pAdMKVvSAyJ0ve9yJnAlkBLBwBt7rc/2k
Ou9GwRbRmO1j0Rnybfv+nUFhY/soZJ4HqdD+YAGwU5SQPpoloF62pGfboocG6nkcmFLl5edF1962
ijtDr7EibwepTeLxm3+A3ycDYv3qc+NtBfnm33FJ6VLcvCQoP+Jeb5dcN9O64m0P+O0Kg45fu3ZG
IsKR4qKUNC6AiKUR5tCBKjMtRP107htzOk3h8sofA1lYTL0qzMwEktnMMdey4L70rh+SaBx+2fJl
TSszo9CAlUvjrcoz6rlXyOvM6QhEYTfhQOATCYz/PZI99Z1YQI7FVMlreVuEMiRhdqNLoP/LyJx2
ma1HDd4NzghVO2A1NKpVMtE4B8hIvdk3LGPdmJuiSKkdVAf9RE68ytD/XkeQe1F+heNgu/RVvUC2
eIcvbA98tnHvjZpavYsyl4Je0AnUPeNWo2Wxn3k9dvIgkiiUuKdP7OwiatOIlKIVQrflV+fo5cY/
ZHS1T3w1V3sVn5o8Zwjmfn2dvc0fEFWwwB7oETOt1Qm5vzTF2FW5JcUZriQQbencVU8xOfpDgwFW
+k2Z/4VLAyQguniuR/McJdyUQ+tfvhl1jODsM81pGg2r9qRcrBHLSq32UZMo7yzbDo/vf/JNdIvY
aCLVxUdYp2bJ2JXayLRLfO0TVbEAi7ktXT5rC3R7JWzE85kNifpi89zC/ZERBPfKNt/pI1KoTmS4
U6yPMn5i9xucjBblUd4uPGlZy/1yjgpmzrBU/8amL1dy8N+iW9+Z8UYYAvF/ETmM9sSKwTH3rg58
0kbaVP8Bzah3xaEQl2vDYeiottYScUmUkLz9xJS+//QkvM2M7ExhLmvuvDXv1a4Y+0cJe4JPq90A
ioLHJTmh1Ak5W2177RXMcqikUihYs7yFUrJbNebk5LVbFLtaiAmSy6Z4xXDYgrsa1zFSXKiIAEvt
eaA5BuRDk7Te5j3BkHdH3di0O5IkbZ4mhqRuAie3fsrK3GasZ5dSXBXit2069tP71yBHCOe+DEyC
6Wltd15cH5a9ARbwT/4MLD7ttmDPoZWXdCqkm7KY9QYIxO99BmQcTnugT/joSs1DTcZyjxX/3BzR
t6meCLoEWcONyNfByy25qN7prqe/rouGc2Sz12esVI4DPyDU2bLkIxZcIPLa67fLPQmBaN0LtcrM
+VJi7hS066yLKHyqfqnErmPqvSBuTPQsvm6FE2ziRx+VH6ZlvI14keeDjpk3UmAnm8f+YN/0HQ+P
fGJzfJfvqLcwIAKQwPXQPUlnEFw8ujvw2E9U7oiY+0YffB2hYwrvOCudtGqzxo2K5AJSPSBplDPJ
x4iuv9RNdYTA2o+ajS+Qo0q0SZPD6BB/vVrpmx9CFkJIESEFlJ//IixjkkUVTbgK3/Q7uyhz7cv+
GTa+8CRAB5OWJBYkXhZRui4VLyGUkP3kG6jPGXanNC6xAoH0E9HJBwyxYhQoYkTIwEPvFGpOBfEB
zfnV2e8EGnjAmzdudkaeLliK3eRxyAEf45Q1mO4XB5yViCZdNIrzeeSImfXzzv3MPvvD9xqxSd/l
pk30TPChmOng/RHSKpGYnpsyytM9DrV5VVPkcki1+arh2+hVKHV1CcJ2CVBLEWL+gxdrgqUvPTJo
oX2v3ztL09ewnIIFpXvsQAKPlvvaXG8nqLhROwPuE4QWhU5yZw/ajbEF5eyKZxsltB+2x8MOyVdo
7DAIh/X0ydNLYGZSmCM6JQwC1kEjrbpG04xlp2d1QGpCJ3Ck1X/vnm2WtEq2lWOr4Q/cQN/Sqous
GkfJEKnnxRK/abOlMcR8YniqCP2IJEjxf03M1oDj01ChwA9ne2N6hbkc8Wab8N6t/86afwHy7xzg
81+4oILiwk4372P2po2jkkAm14BaFOBZqkdKd8LQLnd+p38bqthCxrWMibZQRDe7txQuvDd5bgBz
q6P9HT+7z1ufy7zPnFUUZMBg79vHaz5W/7RVDsg0z5tPqHQu60rAClPPFeP0+5g3yiywhsmCSth5
EHENN2y0+beTZlhdCZ4hmGYDPy100RL4dmmYtfHGfp0sWOHYoEovYCO7dw+H8QaEFGZcw+bkgD17
TT32zv5YWF4gThAyIj4wMqrM6+ONwM4q+W5PMjEV1CVgjZecMxUVaHwX/yJb6L5YBzWG2VhMjWrC
pK/OvD1tbblBvSxWrHPQkJsIw2OCQ25LaJrDFSet+23U/9sSuji0uSA1+CC9KIdtNFr9K44+U7ff
uCF5AskZ+0/5jCcMGl0pOESqlxpB0o1pH5Asl7RO6oDC9XH2ipgfW91sQ/dbxUcOJ21DxjvsSLzp
Z1tY1ECtgQfJ+GjlIC9s/8g/ENq9O58QTWBnlLXVd+7Ec9q6qXPllm9Nkjmjy0GrrE3IMnWCAvTw
oXgS8zirinQH6Fsq9oLEPLIfTv43YfairLF0lbNvLpjV5z7cN2aiPHmbcmvHU6uDTyZ4ksGSm8nB
yflU0YXsYW8EQutENHpDRqvmiNyFMrVOnDo00wW7LoU0fbtemjhXFfwt8mATURgbQM5iQCzCGqI4
omi8GEftWfPVnd62xfcY86Id8uJAWdwM+Y61/3TtavkKNZV58K4pkN9DCIGTooaPxbOgN635Nyru
0swjCdg962Hq8JFvvpQd6vx4NByDudzyQey2xYr08/lbW+2d6fa7SuoP4HJLrThEdyunFaX0Wdw6
AQYos+sNXH/XDB83NT8mtlgcokHFwgFYTGMR7PvvAReTCQgoiFX8ohlAAEY33RiZ+Ejr4s8iAEvB
5bFvhUAb7NlSGjRK/KVomBME+yYmJVz/j/JSgcKatiYGXaN8s4QJgRmpYGq60idn6pHDlIpzrzgm
9QbyO1xmaREpG2n+ytlHw5c9uJhNMJDAiVHskIY1Psjgd67x0CXFkJsEoWIHDskR8/n7gxG8Jv2+
rAZcwIy+6zDKHeYipoqy6aKESoMcswEe6WHjdGr4WZNodLM+3bRGbFszB9FJ+xEY0sBAH/Qx0NbM
OCCqJPsnu3OOUu10xArT7Z3n1Cajn5Gp9JnvSr6VTkguh6RAjam7+imLeUWFCXUUx5e9kOREdhGa
n/nH9KXYzZMCQUBUuuXZ7+jk6HRK09qDTPbmIrhIrLkfJUCk4CGwB/0JJDCBbfLxJYGQwUZULyju
Z/qG//yKAVPNMV1XE7571aRTa324KTN+LbH9cp/E7x0IY+0/wg2oPDvNER8D8O4sWPKj6xvQx1MR
o25fL9FoeTHe2bvmuwu/7YxtXk73VOauJwiRLQ5f9dakIMvT0jsy0sj3ttYJJtjirGUNEpB51+7W
/yIu3NOhAgk80EB5UFoVLKKjJR4Og/E3es62JVP2vKdeJZV2f91UZQsiRwDalVfVuTbx9YyG39RN
8l2tMOlYyKp5uvOwZTvG5YcBT+2KFgIWmgL7VcFAd5H/L0pxNNXQZODrgbI1J2lxcbD85wgtQUt5
UNPnrgGUu8BYSgxZaioMDVdQifFEegIWvzzAyM9GJ/qxwb5Eyt43eRCGBPPPq0ilUhkjO6pkDzt3
qD7UAocQ147OMn8n6sGnzJrZx2LH9DqG+QjrYt7Ov5Qf5CbVoaWQdjJK1XR2XnDcuy9uzPI/FDhw
oJFqni8vv5P1q0By0LLO9szGAc72LZWIVLy5B71Ka4SqkjGzkJabksIRBsVUtG/4aVpIHVZDiyZu
pxPgBbX4FUo7vHcG//ueRIzQtzwiYsds8CuQoKSxtGm1SAKpfIqmMb1MOhJZ1ooiuSHlbHna1WVW
b+UCK1SIehN+bBUh2rCS2mZFJkE9KguaRvtygCQRpLqmE+zC8/Oikdm1p/PAeNongT63Lz2h/Dbt
fjETXDzjfD4EvmGGAk3IeGGNRxPWTJlJriDIRB4lyCQ6P3hx6uFxyMmNcGcbNq8IBk1xE24hiymh
hbUP5b4dRlEZGBGyvUN4riTq/uJrgh6fysxkKw+zeNO3ISzTD0+o92Lka4X1xAQGiebV6mAemO89
Skzq/E1tHyVXXsxjYCaXCbQwyF+J43r40MX0+FRH74hojePf4uDN7TGIaTluH6oNdfEJO/vukUoG
8h6ha4Jl8Y2DWIZbcVgLjUIm+BzVlr6lu0RC0ZR2kItxj8+NjWq8ECS5/19QPsrH/toccVEPbUwY
Np+nNlAAdwlP3d/7/VMSPRQ6X/0pbxgwvBpUXuq7Yy67JQ0k3fYigGJ6HhN6NGdgafueznNwH04t
fbkil45LEgG0I028LkkiUJcZUM7e6UMPJwkqBO9oDIgCe/XXTp3SCHuE0QNsNZCyucVGptASyMS9
OZGUbJyGRozyp6XnZZg+kDf9EGy2LdpsDDQqPpl3QETRdsRVTG/ZuvtEibk47/Vk37kQA19e583d
589s5dMRct84PfduCW/719hOkQyJAD0yoDP8h6r5sxIhho1lkopUjffE+n4tNQGxuOW4u33qxFiP
n6iV7+onkEhmeOkCE6NU/lDqEWldHMNwZYRUGqFDodZ/594F7/iVgFAhh8Na/2DLOqRrc3IaUnOS
xFZjO1K2TUf1CVv1yC8TWkbb9p41rG1bBfH3UlzzLf0XZ2N+aCDFVHu9OS4GH5LADHJA4X4VvL75
6w3w4M99L+kzJjYwI+rpKDjATxlBVg2wV8ZtXQBsTO/EF8HS2styAM2igLsyb+VPsA9+1mYcJkmZ
D6o8gGo3grAa0WvTLr305LZUg2nEgI1+JT6c6+ak3jkcBVsmsAC4k5cNPiUqdLFaGCtcuk47rg0y
5yniGx7snI9DzfWQMKQwYqrLVUtovrcgc6jtSHrCMi2L81qWc34dwlbqKkK+l7uGD+kEsdEq2lqm
kb7tnipnuz4iABf4/HkyXLgtEwtIGqzstjzMKjaVFWnz2QdxJftYc1DTlzqzTGt3lTna/aXad0Vs
cbkePIzrtv1ugIjrBTgaI757yvd6Sqkzb84VgIRztXxMp/wS4AB+KaH02hpvuX8Nwmq4Oxqj+Nd+
/v2TeTbTCZA3E24HeiHbrGCkh9lAM0ok9eLXo0eKrKYFDjv56yHZbcixhSc44pwH/IGQ+Ilssce4
HXxskyj1lStjMtQjyZWbBGSIR6NPBUTI0xIbNm3CjCsaQSILHK5RQ7+oDqLP/y1zn20ZHoCly97Q
HRXo7ctgYzy1BLyMtgMWH29faKX8qbOc17d8+uCDeRFKOmD8WqDkpMvFevePU2Lm5hHXSF1pyYNR
HaumfucehDMk6SeL2zgifpYOik3dETGL+L9CnBwbH0ytXnuh20f9h/qcenkL+g9l6msD4HDAw7+c
ZMD6Ad/MOZ+8PC8GPMqdcoajDKFrSZ1pBmHuK7Jyqm/x44cWHhFkOZ0BJJ4+KNuDWm3ozFp8Tzpl
FZJqQIUi8H/Of9mLu0f45bWqQTHDvZtaPdtMLI/pg9/6Cfzaetru2sC2xGwHMI1YCPGhxJCkPRcQ
bHt0OL/B+oHiWqeIlhVcIX8Q+IYAPap0l/YmVr/zM00FScD6nfawaaFMyUVIujhbew5zkec7hP3f
ukRt3o3jHWg90pfxDK3OczM4qG7J6WbGK3ESnyFOGUOH3fKgSJGnWoYvA+vpjb+lWU0YKlRdo9D1
xA58gK0gpro4ypSbRPlW3xRPs0O9sMiM5AynLBTgHDXzpmO2kam+gNxOMiV7sQQEUTRWw9+wOp6l
lXrWWll96e6w8XvVGT8UHOzqexrfyAfOKoENnZhoh4iZUGEW7n5Nm7Z3+mOBit5dO7XNMzNK2rWl
nxdID0TLnlLKV5nrXXeWxbikxr/xus34aTIwAsgYwGCuh7V8o/tn7HzFotZrqUa2Syqn2MqI9guP
VoFB5ej+q0GIcUIc/bozwpAhMZaQGAULrxIk0IyiDSoIFh+whyyI3/bS+rDYKuD5Z9SocdGfRcMl
4X2uPUwEeemoUdMli5BWEmIkuS6u/WlrL+5juOmalDoILMrQ5FjH1IwT2M8mbBa5gCr6deSJZ2fk
LTowBBltEm+MOf5xECmPm2U4I1JY2IDCJvEOySKR517yt3eVkuxstXm5baVygr419gMOFs1B6iPe
N5gVt6I0IzKMz08meqWhubqeUh9Qp6frOUMuYE9A/dIJv8VUNrCI7QUDnvr0Jci4erMgYdDABESs
etahfTK1cb+tUvzyktByZkZUznLCSWudV6eMiweSOI1z2qb8ymfpde4doCBJbgiwA5D59kc5J8gD
JXa141vVWBAC5uhGIWTcRBfrEZrMNlZSclW71Bcf1Z4U1oAgaxiw3yxo8d+ERjSJidBL8ueKLx7L
D286Hyq6C+tsM4SSuZ7WZdFMqfYdKN8KB7+SjRmj4XXiQMktMjEIg0v7nnYCsyI2lx5SceGdyI2S
6AL9Yny+/WMdbSB9T3K0KuQNzVmUb8G8vWMsqGlrLs6PP76d7uvTmqm7Z4kKt5v0ca/FtAezpQpz
BSqroaMJh/4JohuDA8uAUXjzOB1tP+e/lECmBCjOMiye0GEXfTdkCakaCWGBYwk/KuPyY0F5L2Du
ASO2QCphXfner9xXfRsHaC2B5yeDLDwHDdkMiC3EC4wd5QjPXhIq908779ipRcWlY+ieH97A36Pq
IsOLysM20CJZHHa8fRrxq2Vvqxx9a7zkR5AEy50XAfxLBeAkS6zVj/J856Sc9JncA39cdPi22WHF
kA70KLYX4kUheXreEwJT+eIzQBrzgnJr5WbIRk/NjV70WkxSSyoCBkpcAsd/zq1XsAHFnyOXWxCV
FF1gMH9K7NaNvFO/QmvSOhERTHVFqMv5Z2NthH+EqO2eUPaszJK/2ZGfyL+oxieG4mHgeUfmSOts
1JcBgdqOC228SX2VQPSpTAQlwKNWEfWsQjO80bt/DyDxaX1/j9e5pPK/UU20SiSDqVSBeF7JXd8M
8LnNeyURtLT5DCRJWdF0Qd+upOMmD3VlxB3h5A2HwpuH/kHGWPoaKrLTrRvo5spNXDAq9+Eyf62v
31jxQS20SKv6Fk3Ao7jgOoGn/w9r+XVmHZdAGVg+f/oLJEoZmY7bZNIua6MQR3p9YeBqloF3xyGd
9tblchpM8O1kNzqjZ9E++TShcMXa+1uAdEeb9Odyz0bxRll+UfwJCwHb/ZcuBH5NOadtX+5lZr4h
GultGPxDax3tloO78A5RZegMEibxo/r30ANewJGVWFDJNAo2HVOtscwUKr3DA03chnHKkqjEU5YF
yRJDl2xyGuDmMhFoVl5+6lFqjM+atRh6933gs025iOSRPHqdMQz99tP8nWXTYz6DtwXp761Gy7pg
cVw46T8Bu/ki/8BI4YAlLXPtUo5JmM9r5ZYuEYFYgOkHeB0eiVIaDWpBBT9hq43w/jtI/pPOw43b
KV3Jpu7S/9YIyJPU5GL1vesjf8DItonPKaAE9h2vCxDy2oFaWk4c/iK4ebSiofY4HQTlusxrK2Hc
eENgiZd3HIJUn98vbCYoU/yjWJy1OrsrmcdmZ0nvb6yHSKRRCrJxr+qEJpMg2snovXtx5am4DJCd
zWjYnztF/sD2TfnG+fFZ/SBvm4zIMBXfVukmXX8IbIC2jNHrheHJH8YEnTgxeUzDZCzJ3MNNYyat
UHYN0mJA2jwSC1K9yiLGJAvWhNoNvb3QoaPy/mvRFQNqIeycYlW4S2VWVowyo+t4jbgO1SxmtwjL
BRWuS5vAuMqDRUE4fVHN+nnwNwWkHhJFFsGNC1WIMpFjO1CqytSdHfVeq8lPngTN+OhnLEXD3WEw
FOlY2EANRyT4hGB4EgBQudeTosoTysQIQJ1zLf0RI2BVIbMuCfphmCjdiA9rRnaShRWxZf/+sSRx
waZJqafvSH2HyXhXuih7fNLFloAMWNBehJ0U7EoMRUTXNlpPPh+/nXHThx5WiFy5J9yr8Ve+anRB
uljSictsf6h9Xin8X3EYU3V9H67KE1Q+9tdoKvzpnC4NS9Kv1pSsPrOhxYdNDXjuRpcfsDpPoIY4
mIViuzWO5sZ3Co7qIlpLMdpuMNAl+3YNm0pVmfs3Kh54pU+RrUEsAPVUjTc80gFCJRne8WqzifLB
IsGqI2v3ryhvCIDnb0B8j47mvKP2OJFle/CMOFYQarbzaWNvHy9uaXKdM1Uc5JZXOWtA7+fkKXUH
WxA47z9KAO/hfv1w2XlYH3Km4KEabICwLN4xgCPfSrh3zpGAZoVoRoEgMqr3wgaQ7q9jfVYrXEgO
GsoCEDOn//MbF6/0WlTS/0viDOPsjjRPVTfNQ0Jt1PlNqMChLesLXbNwinSlsWZ4nvE31xWDpexT
FG1dgXGNN1PxFK9QQqNl7dePRV1A/YBfdVqTB4B0xxxfK1lW7UQB3fjFGSjQ3stqQMjsJDF7SSQ/
6JTW8ukHkadEdYMTTbIVrjxbIvOENy5gYFe84/VRw1KigFiVvjmryiAbGWp/agxKZcsTQCe2WUSO
nxWiaCuyYQLYnB3waRzwYmKooByuMxOifIN3KN9X4tQJOjzVFlag+CcmpYxnzwTPiclCxaJY+iXM
gCA7ZictLUshpZrhKwatEpEOOZMMf4KP7GkvfKVPg3qClwA8BFk8pR+zKFYMcelZZShMqrLYq318
Idr8/i88pY0TG8+lXkwhdnZi1XAkmzEFdJ02WyLWDPJLA0u/DdHgKl5X+mI4qiuUAJi7siyT/WTB
XWXpUnY2oqwIja/OjoNW87d3pmaTZvY/e6sGGTgWZBixdDzIVQxBFc614VslnYf/61iz7BdOZRm0
Ixq57Fs+yjqTsWH9FCVYT/4dmrDYwgVaypGy+1nKoHZmHwYdlmxNw4c7JifjQ0dtyQN/mJzGuXQ0
WrvBKyHJ5NKG0dlhx2/7ErcqhaZEajVSEvwAHBVY7cChxn1LFKNxk2VNedCLJufihczCITGaRxgV
HXnsy//4ejPisK+qyNRQ+Ba3Gpl7DDGbSL3PqZZDrGTDgiEqPTY75lPM2jMDRxoQTQYPwXxmzzFI
oAh7R+ddvHmMK43B3+fwIEEMxFgO9QYtjtkTCsj3tp2mEATj1WY8J/N+PY7dLJXM2fnTf+8Vctje
fbOTMyGijb7ph/TYNrYn4gOU2ceD1kxJYjpv2L+khp2glS3yEV2C0QzBuheVLH5w6uFASoZa6PKW
7S5Jh/IFqrWTSRkxSF1qel5w9WWvmd4+ski5CfW8Gstc3Qr3qmFqeVzY3/q91Y/RbfdobFlAWYlV
3LJtknt7SR9ytJ1qDJtQdGvAn5tSOLUUJFO9myn8YkNE1zBIV4k4dxIhtEuyAnJZ1lYwDmy4e7rO
Jbmz71U3xsRjPuaeslzz5+cH8dRWPufW495FWm1pm6n9AFtTXqAvjWMuHJnNeY3+VRLVnxzQuNBo
bH0NVUYDbrEI3h1B6YoAHJDdHxC0/r0tyR4PRnGGWy3pb1s+EgEG+AupEkGJg8DJWLmY7lTwd/br
n/JM8JpHbb5Ha4vPb6wJ527ql6bzR5F4yJc4yxYUPSBMzes7JlHkt//RMKj0Bs0RspYHTR3nlUHo
jM7JDIsHnJb3wVLr7XK4nnKD58oWWb7VJ7ajShWIV7SurKvzzipiF27po95z6Yh7SJK6HICsaNqw
NnfqraPuJRbcX+tTMAzTFjcUijGPY/IyDV98FaTTlBmeUQgj43KsXpNZQ+m5WJw83xY9hCAEVnbr
6Tg331pPsUYurO7La1nF+4QTQ3xicxd1txUweVHnk4ElnefMI6MA4gq7WThi9nLpXkTvrsTxWpke
wkQqPPjJsgu1f+lzDkyurRSOujOdO+j1YhcQ0jmZ9/1Uso0SijwylrW/7o38jmDJzrR8aICpyjZb
+MhLKEvHyItzdb8t5K7mknQkbpAc0uEcsCUDGSd/R5blPtGIfoClWMdbKddwS/Xs7TTntd17nJDQ
Dj+OLFbtu8fco29Xds5buM/LEu561/0vgnK++S9jLqE8wjUzBj8JXt/6NrJwmb+GTVODhuCcLkd+
eC6926eiMVfdMHSIKvKZWGx1jhWvbqc5lKp1Tmx2yYzV/YyZGD5vQfDax04C1Eyk1CSH8f0eIj5L
SPuP79oJyp40oynwWWOYoAsh+yM1VCRIXKWM3e73OUYJ8mvAVQzhpefd1xIfd0MQVqjadIFryJ71
D5SxONj5bMjqw0uyBq7+YlaECbtk4w7N51WpLeGHV/201b8iHrn7Z3lstpjKQa5AEU/Ewcyb/nwZ
kZosM8dugJPfNCCxkB7Accja1jWCOTZCEwdb6bx0pqs85G9PBjh78N80uoKIXZRN61JXyjskrZr5
SYROMcPTzmgw2HwCZ+VMvWWvSgcbByMyL3biHAlNb2diM86ujnmLyv0mim07UlWrA5KsGP9iCRXG
HyV7KO/iSNbVpgwwzgBrjGAzlkvy093Ey3trJm9MSUxu8YFSwpesHzySu2ZFiAkTEQOaUl6AthX3
kWceRc4PBHkK4F2kQAG95HH1TcnHrfwjtnhrxFYsCI7UFRg6GDr9Li239HtZu8zql+C0KDWLL+18
3MYNdrM281qoqirCNuosoKC5jB9Fek8LGsDy1IH3fMmnfuhzpoFLjXjjd/cH14ZHQJUoyLnBDGY7
52rPHPY1N23w87JlXWWh8ADC56ftnd7DpFAcWJ9/L9exj8ctStdS8hwE53J2TrPMoxEgzsyo3l3A
5gb3MMBIGMsOrcTstzEiwxNgF1JzBL9TtkXpOuDxHM+iGTFVLl71sgUljirBsyff6QZf511MuWb3
/nEQWDTdOY2WWr+BDE5wQ3BnqiEzsz/zElELHrn9+aBPZ3b77Raky/vGaV9OsYP56WjcOsa5IhI9
0lHPKhV1DhC+IJA/Igdj3OIN/xNtP3bLGCnZdyOX9C8xZKerWj6bX+wtNZbvv5zvbU+NhZH5vI7z
woTTBuXOPM3J6tcjz4DJMYK517oMAPBdOqMZjAa7Tw7EbmWv6ltLJeACtOAe7zEfE5g/k3j7EUgG
RK43rAVub6fXAKfECD5WN2NenktaP0yFWqQYYIrG3ddHhyT7Emu+QnNjZ4r7WWP3Gh7ndNjl/HTP
6F1NMuSkzV2dPrka5l2uAS3qabVSDPaXs6BOTkownKgh96GTpDeBKRdXsUKnXr8jIgOXFfnY1PAO
x+NMoa2U+Std0U8kdfzdvPdn7UpCr01wnLK4krcigmD47v7WaTad0Hh8tyBGsbnrn8sy7nwLBX3l
F+Lkjeuhja/Z76OX6D5OC91SpqEp6VuyShFOuPcAscAbOj5H1siQ/tQdPUwkd5vSOcYUOhxxqfyk
NlTPOfI4rC2Em5wBDCBfP2EMGWWfbpEkbmk9o/Z7MGAh1bLCVnqaGnRNEnFYKg1oCNDXv4PCV762
CkF9ytiD2oq9F+aBIZO7PI7T/a114pUz5o6v+oZFh9g+2FtCtfIOmtcP/GzGiOND9QMLAyfv/mIk
hkWGfVpWjl0VujCI7MpyKaBfY4+xg8xlBihiOCnj3YweHdOAsCL6OR9JWB75qYdEAJDd59J+KsMi
Gk74EUSQFAzuoULd5rlRXSAGo3AG/3iHKUlmigBWhs2n0yldF3Zr2xV0mCKQuS0hLdqZwJdF3GnX
+PFBoIyFh/RdOXGZGzRd/cKCuA2WRnilr7thJSMUqMQQcHB7FKsN4mD0KTPIwigWW8p2cATxt1yF
XgA1nrGShbnvn0yN3XF18xIc6wJuW8hn6Uu6V5VoEgcmdyD7cpu1w5G8JRVNTja3oiA3o4wMxO+n
u+Ci4XzmB7ibhJ7YtmAorfPgL6OQAjyfbGaiFEDXgmu/ZF61zLIOU2LD9Lx7h1dKAbtNBbm7yqV7
CRhoIh2yp0laYG2QnsgRAKDIRoschBOrAzI3CetKexUR1NahCjHlM7YgENrlx/Y7aYgsquKXtmm5
FZqllr14HH5XEDP6uFbAJ/xr8VEIJV0PXjx+HW5bUSjiUqi3P19+dgc7pEVW1a2jQg9MZhtU+Cy4
2Vs97vpUvx9ds1veLdq4u0OCQj1i3mD+0nwzjXp7oP+gJ/lQ7clOeq4GLFppgiFt7XOZhgo1+cJJ
mMuStupeJ1Ua3+evcvgXW0mvcKTFtJA9a7hvhAIql5zePEPtCM/aqGiJLBQpqLYjQUilSb0+TlP5
C5jBV6XQm8bIT4Iwuyo6VMoOL5rwLpw9nSNIbmRl1Z+U4XuvJeNDyCcXJnwGRaWEpbUI1mcouFdl
oeM5CJNk50Mfy0eiX3Dt0hVuHpmEzYRgqBbaqpMtid66PS1FkFVS6b8KriHs/1FjXAFNUUWaUYP3
25MGE3f7b4Wx62xoQEjOmmypLsG34fOJCYOenC6FTk+oGhviZWVv2LW9bPqszS6PlNHActlp86Cc
Ew9G0TG/vkw0eGBPej5+5rP5aeB6JBTHfETHjMaLLMKaZrEJOSQpViiJGbr6MGc5eCKARZv5uguU
6vJJXASxAHw1TWsMLPZRvpxG+/yWVX6JUODdpuMgDh4YC6/A51dJB9cEv43l0U/BsWMx9eXpBxV8
+fIv6x8quebi01zBShykjlUJWga1L/CbEiuotAH5QhcHY1S8UuPtVR5IheVshhvSfnt9irYLCF2v
fXT+zwF/gvkIAgHi17sFovAZQqngN9Ki5DpnqGPe9L5W6G0jChcr1KnjSXnN/6e+KN954qkrWzBi
Jfp8WZhVYne4NEPCwzxG+I2nY1xdcM+RmOJdprhqOAJNBdaBpHN0EzCkTliJkfapIc6nPH1XD0T3
+NJM3ipUogSyYuHpE9goFIjsUZXoH//o5ecqYZkwQL/znVJLItsIub36QepvUdx5R5fvd2/DLxLS
NNIccenI7OB9yflMJGhUGpOLvRev97OeZaLslSswD2megqr+GA4DriM6aS8wdzS93omrICEd0QWg
OzBTo3B3b61wKQFv2XP3f+nzwyxZiJO/4CFhxP2M81uAoWGFD7jgD/G5lj4xleMdCyN4fKBxzxF2
KRDCRabFPf2YZZVoxBn4C4ltA5F/tRq16OOEnMn5xH7Jq7TQF8TvYngstpS3JWJIjgV42QL8UbiX
WJvDZHZwNYIB69D6IHHdBneO5paQUPmNCj33QU6QolVfsmkcuCbAl7Nmpr5mapWnl6XT/5eiLrSe
KSS+N0tMcwM0DQA9SQgE9fpOFYcoCmn6o2dbQEYt7Cde9cOKU3q+LfMWAxjLw0XImKew9yjcxD0+
z5kttWIrQuqNj911GpJdB4s+PjupS+qbpZH7xUmmfGmJzX2xUqxI4cjvytw/UvZKV6hpT6RJSi5J
9k6+o5tfhHw2Qve5gPcmWmzPs9BwPYkxdJBgit8kcJ+gC3ipCyvBJbPj5J9WyLEnHwuzrai6Ll7D
Va4Ut8gkPo6ytC6918tkt1MjkI24hkP3fjHcJAwxgiG6Wgwx6ADeVtt00JWVGVtsixVnmj/LXaRV
cfmbeVe0BF9QRgaW88tJcs7dyEXNP7cRbn6jU578X3aOjha1NcDaHXImjwOMR8VsEzIeJAcAe0rn
sk4F/acMLUnWtvhKt24+1h8rxwtNDxZwv7VbB8P8OmUoVd0ViszCE6ek8VghkaV/Mq6kqCrbaKCT
0b59Xh06Soe+p9eGQsxFgmDQFWeby4EPmCqXL4yieSCV0FqQVaEsvjZWNNWFsDfgmvCRO1zJpW7j
dupwdrbK/5pHawFfXdeD8YaTJAgKkACZhEdavxt6J7BM0LpczHBugIhGq3ull2VetYLr5rovfUUZ
UnMSAoyDYR++QroVCBkYO34DGzItwar+sNX/ce1DvkJvlUv5Uw9OEatXFlPmw2TnEAdqK//H/XyC
4WO3y9TxC5IEyxwSl0kVDllHV9U0DbAsuxq4A00rtQ6mISTrQV8r7lk7lBANpJwrq3fZI/Gz9NKn
VC/U+gjfdTypqHBsv/UjnajzT909hMBYslcmNVnxFt58W3ZZDJ1QsFnC1Eahr97ZHNuqmo6CbtEd
T/OKT/WOIiW+GgaX0V1G2+OXsqO71nwn+n5o1nyEfeW/+u3k0Ed7capdUPqwTbWinoW03oAg672v
YhMkz2l8ZJ0fmksYoWFSL/+ab1iOot7f0jt+1jYEZtGborasfFesILM/TdG/SH0XEIYNpxWb5WCK
rHjBhzcSGuw6uIWP6Odauf4sCyr8lNqYWkrJ373o6oGLanmrmhBUmbGhgJiaAKlL9zO/n0xLwtVv
bCKx55djOLhnYE/X/T7ffpqkqe+cZ4ZVnQuctNPYXyaoMmi0AeuV+2gYguYqrj02/zI+NySUysvV
eZtDNh8hhe7hmbwac3MRCRsb2UbooH4mWtwnzqTou3TWf1SdTQPQ6rLMRhOOKkfbK2/vqW1pPCD2
vCW3ywHz3owy1eXCarOSm0VHxYOwdoJF/9ka3T3KcZ8Ek/vh3GJ38BgOC/Crggpffdeql+gzNjWY
qAZIqbayRd3o/JF05fvivV8i7SLpnW7biLCWUEigKvRC//wDSkNQ5he1c3JyotZtOGPFgyAuYfeQ
C7OL8LTmRsYhObEs42f219rElFD8uboAH24O6iGECVT9PfO9G7WLhQfO/BNItlU73GY8uf+PxmlU
9rKKJhfFI+I++gZ16kEO27dxR5imez+XPKd0CVcBBVWHcoPwzz5fjFxKYxw1nWWGVf+VcBAkwGNw
vQOcf0CCJf82u/y7Lc0FxPwbxYlPCrfLmkA6sgwjW6L6nCwKmocpY7OKfTEguFNKx9djeNY8a7GU
MmA/1O4bHHTOiyFjeL7En/licqZIwvbQ3kFI/6/DbDP2YcGejCw06YzdAuJENPzEXcqUH88YQDWb
GuqXifUabsR5MS/Pvlzi0OxoY2rwftQ/SFMHdU47n1cx8Dfcsmh+73tgxIuuEM7iOoKy55P8IlSA
Pv/WiBZmMpdIQn0WHXQF7ox7zlD6xaFzKDXHVGnW+8MJdUbatrrKWNsLy8DHMCoHEgMr4cFjIxFU
pA0rG3OnDiU5Gn5zgPXzXyHr2w94jIEl2OXI+YB4ueFe22ZNPIuNlf+81w2UFxss5YsgoIjeODE2
KSuhML/zi+bLIu3rRmbO3hExk+kiT7dzC/wigRozLqnokQCqRSo4uvbkE0tIfYVR455RgBUFPsz6
9HZOHqBZgoPI0/Yu51VidOf/qQWiLgveeHA/Bix6HOWR1uymugN6tdeXcnzh9CWDECggJU18zCJ2
ixc7mCkaZNebdLWqqMLvlHMnFKTLB7MzQNHGGfl50qQ/tZwx1THCvyHGu6QdgnRTbs38Ksv480ad
CaQ17TaBz3l/H/cMfoYP/YD63i5mdBmB6G9fxqqydn5m5KGNLa/clS6NpeCnyqWC0b3Jw0w/dEpO
F7XUnfcVxhR0sM4xG/cVbd5oWSgLDfD+xrSGkuY0qJZFhCIfSX+AQeKuc/fPWomBFWiddyE9htQy
A/LZDJ0j+53YXJ7+Bl1XBp4d+9QcPyLEhqeELsA3e0yyqZBwGG6z6pS33LRAWhDam0SHpIjBwRZf
H3NW3LWQJ6nk6DwtY3JYAJ0oncWJnj7NZoHjA5F+5oP1K1z0Zjqyfj+f7BjogNVIO2eB+mF/VKZb
jALWUako02vqwVS/PgQoC8hEA1/aJmcbNdGvgKMglbotapta9kVZQfhfFIK+xMjxooVkqAyIPecW
r66AkVyZj880tDqgXs+DRd3eZJaGGbryG8s7cNzdBOFO1SlFvqr4me1TZzTC97jSoYOlOBun2iQN
oXMwnnq8CIEWshVsFsv0XKQ9PZ18/TQRA6wrrrxdpDx7eIB4GyY2Uu1rT82sm+qJW+i8jbGwrVi2
7/YaEwNUrdjMPa0/AD4xhoqNwsvOLL2I2brjBH4wr6NqSXQ5uxoMrafpONK3HSWBd0kM/zH5gF1/
3kadgHeZuKihYA3TYkdL/xvE5OyQOio2/YMB4nNz++Qr+DGT5iIicTfwqOHz7nN++7rKAPV064ce
5bsPOgx6rF3glqQlr+Y7XXleIwgWzRSmIyqjnzZGV2zGjIaqMfWhV2u8OzBtZze+xq/gcKdFEbtb
l0q/RQzzbLPgaSnmVXJs8HbK5ooeMPQRHzm3SQQxeFKpnmMs/xOuo8RWyJBjG6yqnn6hV98rxOi9
vQgfX90xoOKUKoObq+eltJjbq3LkiReDWRFKKeKOAjqFVx74wrdk1G9qo9JyQg4bHr27FjCpY8WZ
7s08GecVMOFf2iCuvB+pb+Em6GxXYFsgZ+JgKjUuY/T2G+hN8mGaLagR9RyN00Z6I8W+cabVnwe2
422Ms/Y75dayXNKu1z61TJ8z/OxknX37/9swdaycT2mX/MdM0IfivS5+wXqlPl81VD3ZPWJU/fHP
0E2APzZlNEFLgtR/Lyvof1KVsmYaJoOGQwz0eju5T9NdgQmU/xQ+hzOR6oa6EdHrK5pBISAMzFYE
GjhEUS6siz27uENeWvyQ8WOMYgcy7ZbF0Uy3PoGyHJUp/uyJnCIhnPQ5OQ1jTcR8nbxo+mPrUbhx
M6J9je32TIYN+tLXGs9gFyc6InUiDUsWOg75tIBEgZtz7lwJx5xMf3Vi8czZmo5HU4jWcB1bCcxA
Y9utetL33sTVZKXBzumD1pf/8869nJMmGIWQcXSERJHlBNZC86kwT72CiX34c1kGHKg2/xVXIo1v
Sp+6t1c2JjNnmBqR/wKFqPAXeM8Pyae71KPyR9Rla6ApIehEzDqa2YnpKAkOldLiV2iBsZlC6NPe
fsWfjFAALk6AOJ205s/0IwAZR8e/8gOPTi8gwLFDOECh98EMxjV9Vrn4arweNwbBMgCutmh+x1WE
DWDLmbJG7H7MnhA8E8V0SjdHzl7g2Kn+ZZ/cQgrggoQpXpLetjxKSIadQ8jC2H7WOJe5b8PTjpQD
QXk11x0A7RDJgnGxkU5f/9OrmkzzCqNCaCcMFGcDd1D2HKeEx3o9TXGF6yiwiyIcHCUDY+91n7TD
W6VQgd/Jjh4TTNa5jLaB4sGfHtWtunUmSeIsBUoW+PUlRn6jnuCy3SmNy+S/jX7c1o01DYsHtTH5
eEFGx8wA9oNQj9i/CXYmx7FlPjCqbWo/R+77+HQO/uLHsgcttK/Xdh+Z1hgucmLXuFIPLaRT5QY6
oAAl0tpDbdyfQuexEdSd3sJgVBVWJoZQuUwSQW6wSRnXbMLSgUqhOziBFiSOruq0xLI1eHMcnYMg
ZX2zGlRMiPbY40oL+JReVD6xxvDX276dkMab/BFRy0zAvVQ0J1/5VxpUSVxKlLyrmOvlRorrRRPr
xbUCguBoveQ7HxfJdqurRT3ZENx99imxP3muYT/p65eXz49xMJqN/S1pYMFslR4oeur0LUqkIUZF
eo5vkH0978OMZh7mXo81rXVFIkEH/msTBjhNmpuSQhsRKSe7bQXBQNcuewheaDe2hgsOa2WGTXJG
p3PbmotR50lMSejvRa2X1XX+qEq5nINsk3g+gsn7h+uWL+R6Sbo73FuQ0BC4A7CXe4yhboa0ncv1
z2Jv0k2xysaXTGkhmgrQ4MQA5K2MtMVsagJrnWE6/z+XkoVqOQ9fIBy49bmI8HRWxD7MhSDoWyWK
lE0yP3qG9uytt0+WJH3AMutQxX6eEEO77ZDSlDAJemQXSkq63FPkV84fH1/nhVMLpL13RYIkiJbT
T8RJ3VQizxJY8ZTAxblvtHRZZnQRGItA/K6pB6QMkMg1zzCtZANXrgmI+EvEkcxYCXUMuGRYsFsd
De+w0tlaXklYgCir7ZTo5c3lr84/ibwL0i0idrFz2EAU6GQST3XYozKXgrfSh6FzRzCCVt5Tktj9
qHdGm56GDsGUlzS0t+qpgzjlcpmTUK6SadpTSQwBmaNOEfTJiIUodUq4iSVR9mU7Z6DxnlvB3dcy
7BdODKArtp1bcNAgIOGmR582EicJAuHoCos7iq5KVUtwV92xKm2xQdv4/CxoS7fx5w5ojTCBqD6k
SRaKuhJcKWQ+AFTQjLAJd5s+n3sYMUs/qZfaibNyluENf4+THGKIjKMPtp9izLlSnITZP2Qw8g9l
6hXt+eP7PWq5a1EGFvxYAEK7tKmDac7c8up+Oqfm4HFmDPeZI+k0NopI+JuotqqmVHDJqFxTffi4
Xaja8zPTIXM/NN9LWBS/jo2E3AYXjToVKwa2BKhCdJ0CptGoDi4/4Hx3OlikRsiOYMxGLTeNSYF7
pliOWi6E7al1SA/78meqtSLjtHyE5dkxAyxSCL4tJ6LZscmsCcN5INbfsQ/7Bz/0F/dKnF1fQNeI
BCuY8S+yYHQ3lUOoa7nsynYOHgZnYEBUWwm3olsEaWy3ItCRuzSelTXsAG4ZmoOpV9YBJ/TGEPPN
yTvaMrZXo6bgkScs5zlDpq+zocQXEWVrGuldYFI3/4AMYxwRja9nDcBmNQKCXCZj1DS0Sg22KwI6
DG8ovmaRqa6ZofN11RsGmNdX7X24FKcFRpcvKubyYJ3mrabVJHUwAGfFWkWyDsPfxoxP+JHb++Bl
khH6cGWokwrahtv7OUN4X1ngMLsK5vXBLG6G1aQ/n21sWKtWjIQIVOW9OffRVLwlmHvw19VYwOmU
qYm9gUPbLD/qGISWXNTw12Eot4pmkQnAs+gwRWgX8ZULbjklwlS/czwgv2NuFiJ0IPmyNMUTN/Vh
Gp6vpXTv5p8HaC3U+9c9Hev9eoDvX+/eMJhpyUaBTUr19xXbDTkK6GBncDbaD2/mwhc7xSs9RXs4
I+TrkXrfpWA+6oYrp1OMKMKhmHd1Aewsy79zXCVDvQzeOYIUMZvP4pV+jRr2gAl1jAbO5YxMSLyf
TmiWuLMxRsKBu6rZB0XRqcIHRYBKkOzrL7+PKlK6JlNkDl+5tEy8t/yNIWFZh8yfWGeR2bp7P/DW
BDyznw4oQ3E3tcC3qxIYA7/ecH7+4qEiMnWkOAJTSg1t9b2j89539aqddQVzjCDtMwWjnlLe7VR0
T5hkZjEkW5eaQU99wfI17tJ7jpPbPm6NAcfsR2KiqIpzBh2rjNi3z2ZwbhsxOYKQbfJlDBEfwOGZ
zzR4ONQWnSA7oP7MIvkGqiWrhmQmGA6y8YuJxSgeVQq3qr8TTLvZKPEXkjGnEj9aZREa+sVv+2MG
tz4kR3o/mftEueRogMwIHmFrSlJMnxIKCGOUIS9vmItz9iSIfvyR+VkEwDrJSnl+s2TxpYq4016V
bCA8r1nkQxBUIn6Z1m8DC0AM034ETx13bVAY2hrpRPGNWAE93iFAA6VqiMW2BRhVx3T5z+HbT1X0
HcwFtAD9CYP+d6SAnWcVG1r5822GksxN4vhgRUMmgok/LTD3hO/q35nh34PB9U1XRS3tnbkIZYQ4
HT2dXI/pGwbpBNOKcB2feVBbYRmQcPF4w2UnjILcBeOPYzpHLm/CQo/gEzUo2nOxkk9yyo1TgoDN
8TMtIjbC6bthyALdL7ok9aDwkBuoPXRZtCLopIcSgLYx33Z9JXRUkOyXf8pUE1gJhjgRuct7i8Gc
qAr9fBhCd2k8Ljw1ucd0a6SxQRBoc7lYJLgzG2LxJVmprM6B7MgGjiky4TyZV3aRRLfOJt9r2CiX
1Vz0NRxwHE6WioyfEgI3gtCHfoap7c5gf9FrF4ZqdxqBP6xZq6wiakp6oHCyLXQOOfIoNPp/H1JX
9QwH28IqB2H7ikVRzqF0Sr3sk07YykNz+GaD1T2cm4EnZ9okhgrpRviPqu+k0oedcZ1idMvsscGU
wC9ilyF3PpwMQBX43xYIt6YJ73yIaaVrDg+ryhwfH16Q7e4q+jlf5cTwElppqGZkoaQmLC7RF6Hu
+VSl0zxqHBG8vBuNDzycrwKaW7xTy+53fQ+n6gPTLOJ3GuNis5w68gU6lAArJSfx5Cpc4slATswO
bfOilCF2VPLWTloUdgSy7Fbx8++lMv8dEWX9hAUyRIl6CTlRNNmZzDkt1aMgS8TzU8dK0J6DODel
2/OPQee1kxInQ5ngkB90hGQfmcKjbQ7JkOGNySA42LIIJZBPz2PWfwAWl0bg3mR7PRN3Tyo1LaR8
qDDuyldrXGWhwE2J9xOVwEjwzzdQ9tfCDiJS04mtnIKRH19Qc2yZyPDSAdbbt8k3NwHVrI8Kh5eM
/yk7hCfCqG3EV6Gr50af6NiDGl0M7LBTXjtD/zinGkcm5TfLhqOVCotaX50AHwkMd8gfAp3wxVh+
8ZURNzwMX4sRXOjfzrHHmjvgqzkJsF7lVIj3ZxZRdzUh9JyvaTEsJfCRfam24fgYbApIPQy1LQe6
wpFpNSuFiyN9buPpOOdKho0pgx/i2m/uBFs3kutEcJq8OAitUUqxq/g4sU3+h0VxOWEQV3CMQWIr
0PPzbKOLpO5V574xoJWFP09OF3vgPVKzLkKQogw0MNW4FA4DuH8bq6c/3FyVeZTP4WP0HCvQ2La5
Al1PznRVKKevHF8Y29+uzAfBYkSgZRHfIcb3DbgeZNpcY0rBldT8jgLPg+NRJvysktJtUfi1CXVW
xaWWIVvMluKgj4pjOMjqbogm+j1ajY3TH38/Bj5LYLZ3XjmfaDfZ32pFaE/pX3YCJmIKRlJC/FSC
1E433tZL6NLj89bNIGqhHE+Mv7bwTAlgxb93oCzL59Y+PB7PTIXHsoeVDsC5YEvvfgeSM5n2pFez
XJSXwq/z5gd2C/EGU1BOInj99/7qtRq4BkFBZCMNKD6k3sGK8YOGtzHl7Je5BqoyztynnAmrz7IC
PwBuXCjj8sRd6ZKoBZ87l2TJ+PW9rFJqHwu+7GovJ+CR4QfwgtumTszamoEOvDMciGn39fLDSKTU
RN40OlrK2nkBXsIKcdgeXmY03yxTXLN6gIYqnxxLl+GVo2ebl6xlCZ0fUjmfkbag3vxEwPCVEpw5
L3SNJ22AzGzzxXV5vc960RWpoCfsM7/sSEZ5DETBlu3ocHOxyE4S+PtWyoqM9laiU52tV6P/uMPg
oK7iXiyecrSKJrRESPx+7/RhMqwr7stYFVgHSQUzu0qtdu1SVY8RDWr+QV6KiqMpNO5ZKbVd2Z+V
Q4+d95Ih8oQEhOw5gXksCKWYFxahcto8VpDjYUB/nBd7+C8SNIjKj8TRUfKn2OJsFMtBJv1j1MDV
cdf+B1PK28iBi83oLHzC176+Nd74AXL1sMDMcdWsSBw282Hzwv8CTneEKOI6rMNPDe9RUl75sPhg
X3+JoAEwfgWI9EF+9NIJH6vuWTwNPiShyGlBK8Wx5C4qErMc+WPGMo6GUvIhSpHFQWR8o6NFtSk7
DflGJwvDa6hT14mn9ZDXbLG13YbLUDBEdrcbhQhbEBU9hLdi4/OpMi0+myk8PDXG7avnH6H+uTev
5SDPxETDBgZDqwlEGrcf+lil8dcs7NEZLKxIiLhbmoKvE/DR2I4Gp0zcDJ16aeqMDVwMs+nDJPVQ
0p7ebHUE1vUOMxaT6oJy+1gxnDPg8Nn9CNPJfkNSx81rYlN6kYyGVIHEIz18dlzdsl+p0FJ75Tp7
tMAflNRF43ER3f3yD9SmiV+9BWOutUzgcrzr7SprzgM9GqevFOQ7MLc3XSfhX8akAJdyTj050Fzy
TUOcLQv2PsN+ATAf/AzY2NSqCr0uq9k/OovUTY149vXV4gJ7ztxQ5AOsoGxGCfShFVnbTOYghGrb
fgqaU7i2rbTWkyPKLdrxJKxnn4Wj4MF9JZJGUgZLexVvnMktaNclWben/DpNTI5hhXkHYSeL0OeA
XHm79zYdAFcjysnNF4+RvXTTDXNCo2PdL2OAOhliwYBby12ANZY5+x5ap9bJjPluhKHfiQSZv8xA
u7O4Tzt/j7rfWMZRm7csGx38wP4sjFB/Oo3+QQ44TzWpQlOMJUIHNGb0hUhJS+UrgR7US8cfkU72
2eO4NmzE9iB7/xxDVYgeI1stGaJ7kyLLLR0aV90rN4UerycqNPvWq8QSiNwIS83J815EqCptpwVu
G7yTzBr+gcq+DYdsxT8ynDNS334mNsuuohQIvGq7Zh0Kf7UxJtwR/NnlmY7hGR9NMAJu2+u7MGIF
7x3uHw5jyCHNvHJPOfQ6NnLrLPC1oOGVMrKjlngyeziezVv12A7H0oQjGT8J2GQztgkCbMs5kNSY
YYH8RmkRvaGBNtpN9gOt5tUtSixQCchSYlio4POdPNamvV43owPvaPlVcSKj2QV+uwFqq7GOt8QW
u5E7hlaWXM+yWgclRl/Zk9Dt/tgaywKTQE4Jc0xWvRXZhk4oHt9qhsvQGWhuhwuoBmix+GiDhn1V
wq4KV3C+TQ/NV7QKUbVHlQP682o1jN+yHLxAJYQZK3zMLbMBggz4xO4kCPSGLcD8x8YZG9KK3yks
HLFRurU4BXsREKnmeYwy872sSDJuKqqNgwZVyHmlUX3i8hZ9Bn6/yhc5ccYTdCpcIKkOp3TNKJfd
gYXQk4Fi/fgYBWVmt1syXJYm5nb9zXWm/5DiIgNhfde2IG9kqGCXKMBNXR/xVFBucDFtNvZHAZwb
D6nzlxz/50mH13O8FeIBdA+AD4+AWcGx2xV0T7M5tW3RSlHUC13ZxxBehoxo8fCtTW2TAlQ+OaQj
g4Wxfdrp+lfSh0VhOZlnNbiwOQXrSOXXUuh4l9REM2FI/k35AWjHaNLBA03BdRi8M3sPoIJjqAnY
LE/5r1VvlMYJ1HCtxsOXgFuhplWkcd86U0+vq3i9dWtqtA81hWL7t6/FU0bRCHLJ45q9DcNhl82r
3pFuDfZfdYvIp7PfmAVjx5Qs9nK7qZo+WRQcswfhw78gsB+ZPKk5YmNoyS7lwK5K0oggfiYYZs7I
y7tq5Mys/lrydfyNu4655NrmXxNBByv6of3rjlcpZ0gjVm741OJfTRRn+QKu4GOp+8QWlv26n3aI
8iwWsGMdUX8okrJ+84+pg7r0LtTFrazOpxYVrfSoEP//dDYptjWAkDSwQrR4chVA0dAQQi23JGez
VujI96JbE89v/m3o0qcHsZkeKHlWzgJUvPjWURDOHRTKW6jjgr38BTtlfwaJEYgVvfRP9R6Auw59
c8t/ElQkcSXn7RYJMcKVGYvwybH8RwCPnluB0tPqFXvJGhxgWp1/7Izd2TzMsn1JCPBCV2L7Fb2M
X37j9qZ51rz3GGaXyZ6jf6cfgVuCrwKI8EWo2d3QRI7zZ1sm3G7zQZDwXYGuEUNbMdfrvHmd7trH
fjmOcT+zvGtH8Df4rd4dmI5cif48X4eZ97jMwi4JOnOsNABdVOTdH7NAaXsrXerMeUAJ9Fwne2eu
Z+Czjd/9DyMWGX322dWPMINfACyTUNm0pBRI1xlbv9FsqOcLzEe1NoVxA9StkV9EzULgB3fPnnRj
CSLbEc9BJpHaHzFuDEFdwnjBsyWT/mRTqzwxPHdVmIrqAgPDJHHzehnTD0Jlynq4kJ21gFwXhRqH
Ueyhys9D6byDIYbEAVsOrh0SXHaCNm5kfAn/hFYZWe6hMsMY0f5yFbChXXsPwVZRSZrHm31Y98om
UkUBMLGnBUSpUz0aJcAXWgU9a9XOF/tsur01gv+SmpQz8hCEnU0PIyFfHo2cFNpR8qkq4Ng1KD+i
wxgN7jhdsoXH3TKjZt1UavXuX6rwLDT6/rMgCeSE0EaMXJJ9Q9VAS9lyG4+QOJWkE4e/8+jEGxrM
kExwvxv9JWkX7MB0fQ4DqA0+dW2Ifgu4LIQ4fktj84w6dF7W5Xd8Gi7sM9GCV87mQ7fO+SFjTPMM
PvU4874pIPa0nza578zufEE6WQbUQ9L97m5aAHzFPTWg2Xwhwa9/sIFKpmYqJ7l+A7bQoGhhSw5j
q+OjVzxr+cWi1ln4aGzoGBieqQbpsBatNUhgK5K4m192oIsDqTeIJ+FD61Gd/7aQVHVbVI47ujbX
SdDsuAWimBqnmR3tQZEodkmJr5u8FYybto1TcgnqbXssQdq1ZYUu3KdLnIJtU664T64C0JZAxfg0
LPBFgRKZgn6JeyFea6ZSQAgzAGpunwcwKYK8XhTFgSaIrkXeSnbVZNiXzHvbAjqAiX4+s9zPFpoe
FAZfEYW5+YfwC3lsikp/1pPnL5UKlQux2vvfpMNrAuhgEH/R/72injbZJzs8QsuMD3JDwXvJxGqo
fo0f5yrlymywVs7koagQuiySp2srmmYC0HUc1+xmTX2C0pecpoU99W8iFU6S7eLdnDXhklYVjs7I
Jh2pMlsYGn9px66Ny+8Am8i19XB+/QQCiRNPRmqG8/Pkuq4kKLNk4lNbQxiSaU1GbkVLHjnfdjCr
eKbvuOWbmA78vHo74XccYXXyrSZqAXNWkHOA9B4L5aRZ31c4nqHaCL1mAwvG1iCKGyGs4nZ8qtot
SQmuzDGnD7l+/0iSFkrzZKSBA53I76Rcb351tJDS5DpMd309inc4pDjRnSDcL3xjhISluwPuHfHs
HYxMqdFHFbnVOFmCmjxaYLsexB4kHhIvWPUZVfmbzjDnxQ/JQzKLZcjl7MT21xhPjg/1hcxQmBAE
OInqS6O0rgbG1+xf0dG8jAAQyYxIFG6ou+iV/lLqhBvG46eck3VCQ+V3rg/bTVSsNhmHpFxqmLpW
FviWpB6kI2K/VaM3InKSZmDYL0fbEx02pFRxtmq1a/Jld7/6XMBymey9gvuJbZKDgdZoxfSZjoKq
604BM/VXllzKiCgaaZW3mQ8weP/EteEA7exX5UA4dKD/2fEG5RjD+5F6WOQFoP5/vQkQz62KzuXS
L3ONno3/qaDSq5p81UxKALy4TCDhmob0f9VuEKFW1TlvoMoWF5rt5zrfOFdpzI9/pd7LE/hgO27D
+fgU7WLRvEpb95iL0Z9+ZKVQi08liV5rKbBabnVduUQk6Ck0osV8JviD21Y9GH5PTnS++2n6mre1
7CQkXGfK0euLxmsKQyCd5E4LXh5e0DOa59OJOhznKv5U1nF7hHCpgxkBH9V1qUvNFeTVlJ5wj+Rl
DEq3nEhp0xZagDJi1i+x1kH4hlLxfiI5JlsnpvNasdiU7Kni2OqKWVBe6AOVSv4gnO2+4FiXnJrG
KQwdZ49+V5/sDamMezMreMTyEPduCOp8Fjk3t9d8STcJiAbgPFbWpZ3kTigP9gkK8nUC8kt7BPSL
DFWjYL5Q/yAftdBYAd9PPPCGmV4OW4lpNxiGYofiVoau97iQS5zl23+CPeyvaQ1gt/G/u96ZMqx7
i6EtC1zTiyf22nkQOnqARjlWy5NySxrMMWORPkjNAX2WZ++pv7A5PzBGs4za2+99CnaJ6jVPpIEE
D72YWvLPqoqvnM3k53AQaqwLNGWnlVkvWnRhVsfK+txl4XxI10sX6zceTf5AofG1VBsR8+Hth5IM
Y0RcMWQZ2XlkTDo2tTtzUJNDjzH4aP66lZwL1U2N5uDZj7mZppT5Ze+mgOanMsuLNbJOEuD3AqyU
Oi2YdloPgJ9w3i5Kw9URNoH83RxTpTJG92snzRd+0JGKF+leNP8s9qjx+btJgcJYkPkJ64Z2pfhm
+PxvnL6Mnkc0Omed4wDnqI9hmjI4eVmLChJ9rwGt5TesBFv02vaaeWJ6AtntZgA7pRQdOVxBB8NW
lITBeF1cqs9OA9m1JitVCU5gzknd1u+3swPMoIlJhqJM3o7nstc2H88rHZ1f84R0zdQFFmom4Vc9
t10cejDPx86IKbIQmphJjg4HdU2+6U8u4QpDM1vrZUk1hlPzv1hgaLfvuiScstAnYS5Hm7ow9Uwy
r11gXeNVPgq6A8YeTLVY0jEtd2rzJ0746NoyKDiS5Nwqf3PbZd4AnPruSAU7oBs94WQOIckCyyxx
XF4xi4/8fB7ion3UUzA1gVI75FMVohdZ0h30jsnPvKZwBz6WaOE1D3Eg+WYWwNv9fnJGaY/0tvzy
sSLiBfMxuOom3auVsTCyHFH3SD1Lz9XEobQol0o+ClTxcSfBxln47RRjiFk6EobK0NcENJwbXJwE
YcKHam14drkC666y5rAM3JGNHwAd55jp95qetIHKUcTgvAxfCh2H62w/lSkaP1fWsHje+0WbAEtp
tW2tOgKqMkwarxkERbTIHKX/La6Galz0QzfCbCMPWbu9G8YbBRKMP2kpi9PW2DOtr74qHCNIbwSS
w62zlq0Yarktt85CKraRKzC3ySsuScyijfDdnryJNbvbx/U8frqJmqmQ1q51zu9ERqjveyXlYgM4
4A03gz+iKf+VVUBy1Li60K4pBGYtWlSMMiFJkNqd2Y/38Db7QeS/hdN+uG+1r6e9gk5sVTcj2uzO
hFXrGdyQK21rMbXkbPKPuWSVQ2wrvHvfnzYroEDVXOKlhZ2QUjbBQ9/5J5j6KDIgphI+z4oiWhl+
GmMJct/WfiDbmhpQ5d/CHGrDq/7UmJfR1g0XCdi3fHvx9BJ1sn4UBN4gRmrqDs5Nyr4fxTjABjJ7
mM4d0iy8AlUSoTYVJk3uFdH/XvzqqhCmr0jKp5LANaTv5r7B93JtvN9+J9RXXLFVy6LWIghTovGL
q8/St18FHe0Ngx6qF4qZ+GcbroCsTPRlQMyPmEHlXiftR69WUFURbwaPO//zKeQLpYLFJBrlSL9q
FH56V+2u88gwjjsCTJLzUWIMFx1qIoH12iucVbKoJyvWI6ypuZGURaiT6L90I3ZJU0qll/BGDAGT
aA3vKN1vllmsFdRKHtNqLCnpWtSWGcZa0ejM9dvpwCU4lV8r0C9rtfOtgV6qKSiweHjimcoj4E34
yO7qaCaK+3MWPd9jJl5lrcUmEKdLiulyNKnxNr6JCAG94zPASUhAnJPDWpkb1BrZrBDLxJofbleH
2HFDwSopcpmEqsJjc+j1chj9NIyFWVoYY6WDsmm4fmIEgy0etx1yY3ejjuveag+SKA6hTmoKdIuP
uQJvF9pjOHzuJ8bz6YZ2n3vP8y7vGayiuleReiLWqO3m4+lYj+gQ8cyhrOlArOrSxQZ3f0UhhGrY
NV9y2YSQpebr8/6KVvweQhK/AFQWp9aZb1bFORKNBAWLX1xOJ2p0V32ow8nHqP3EkvhB7VSK4JbJ
VndVzee7KaOA9z83VGS3Wg3MNIRpDPs2yZkvJqtffvg9/tFpYThnJ6LHktL5QDWwmo4xoOSbC1MS
G8SZQmlhYs8DoN7E2uBK4JDNCcQ0+9h9UONxQYYUuydW8lLd33tVeAy1nGa2FKcTdnJiq7E4cm1J
RURODLPsrd14zd67Db8R7VL1tHLa0E8LAR4n5O8m3obBhBzviyNgrMD4FmrTQj6Mu40+W+1Yp3of
VCbVfuo/JfIvBD8viLMijXWimkrHsUxUZxurRB8Z0onhT6UJuhj0ouG+j5+pNCxhOaVP1bc9p5Ry
sUjkjCswA6EwR37o83NurZHMRoD4cU951E3TSlJHeFkovp7JI6GPOlfwxWLDcVCmE6H45rvxsjpp
rgcn2lWV7w+Bp7vjNQTb5ic515Qv1SIHjPeK66frW2RZhesh8vYUeeL31bpYAcHeRnPN61auyIDz
fdNGIsk/QYam/2y0nIVvV6CKtJBAlDMHuhoLKzw1ETz7S0l69lG4GKx6yWmwFSp7q16U0QTdaUg3
W+GzubCpB7FWJCsz/gM9RJYZeHCFY+p/rNys7uLxtbhT3TeVKNqT5B0vC/qgt3ZvnEwn3Zn9rDNb
uu+6d9lkjGnbqv2j3R6IGhCua2Y534qw/bxHlrECnjHQMHb8F1DqtgoyjCYPHv+Ln4wnmE3kiFpX
OIc5PTkgwca2miIBnK+qa3f7F8WPKyc1jkVQ1z2hFgtV/Q8ammkXzThzSqOp/Sl72oZYla46V/2/
jezFaKJB1HL/A7aenlFgwNWn1dq5D0ru1Sfz2az16L3wB/4nm3ekepVheIpwY/Nicid3GlOrcbjn
Y0tDTLJMSzbgEXE49HNGR+3my2q6bMeZyjgDklV/VivIojLAdvOpbetTiCgzHH47kEcawCj8y2Ao
f4O3tQLD2szXgbMVGQOpccn1Cc9tB+OPvygWrEQnwVxPHFPABopxaeGu8y/GWsY5lQKRX4QXYONQ
WU0zuXRuVqXNOQwtE3SW6tSjwj4mTbjMMmFV6VaL/lcHVAOe0C8/VyCA3ncYlFRrSRkKn78+5Iy8
ZZRTHzcQG7SAXG5rfR4Rp/i0wf3Ish+uKXCDZcU3OVFEhQcbra2zazDrVfCahRztPbZQX7XPLse1
0+rZnuUrLwXSD1/Q46tooScDiZp5eNGY8oaR87/TfgATmKxzuR6du0YtwwfKXtFgmvelulo8fEqw
vTG0BiVrNPwFcoUz+ms8d3cZX6zkZLPLl8HYavSqk3SGw4p2SGzt/oZZZYaX19hZtCCwhV/tqxqz
ACaxgkFPIm9w4itExJhQGhT3ShPv2H4J0Y1fAlyVXhHU2t4IKGZavzlzPMVrBt+NWSv7lDTAwSmK
EltTSRWtLcKmro7UzMaNagiOtNcPTb0V+etr6tJkLSxLZvd1vsBCKwof2imvoR9Z5dZ1BDD4zOeh
7rlDCB8NdgtnWlIQkUjf+RcLoS0+t2l0YN3cedZZ1ijFxPixt8BVM5K1SFJ4lfEmx1bAkwAwhDI2
7ksvBem6P9yb8kZ1fowJB0l22klFjIHleP8LXdi5nD2M38p5OIHLgb72W3VdWipRgeeYAI98FTp6
Pnq9ArEjtxcJRLA7NESdK8f1ZI2wihIbJuw+HgpBpoq2wGeF+aT54mThGfcSZUUIfXMyN+vwfm8R
GXSZWy/FnCXFnOeWIy6+gnNZf4GexiZe1VPflJbj5QRi8ak8WyqKlsSLQWihSpNSJE2VhnZeLTvy
Qjo4UH1HV7HFW3As9JdHA7gklTvjnBj7JVTpmXaatcAzTDzafFr/frVxDUp6kKwfeyHUJ4Lexq77
I8f2PodlrPVFw/gc80RJshJt+BlnP20ceWSO48vhtnsFZf7lWZMUsgvw8qybhirPe4UgansRLPW7
N/bjrBBjAA2Kd+RT7OztP2sCEuHkv6Rt8nSm6tDijxSy4CNnpwECB021btCyW7Tj5k+BOlfhdzih
gf2YZMMefRUAtcomXrHoPdEFGajnpnUCqUd66UFn2DNaSzRtSU35qsn2bwx2bZPvpP9Pu5tF7ep/
e997SaV2Dbt1osED1DxfvjvX0Pto4njhENsvRx5kCUeFgZZeiCUbtNmZxL9UWBK+OWLs5uHSy4iu
0bTqhqSVh0hxI/hCIM2n3xfGiabaWsvcjck3+IQ+OjkERVEaHYiCVCObjFn6XeQZFiYnlpNMw/+2
BTSQd4aqRIVuvQ2FzrO1TAQS6FN0uideHu2xgXbKFM4CeuBMhGo1Vv47eFrDRcI7hZv0Gwn4yoYd
/lxjTgkvVI+eJPGvG5TqJ9xpgPvdD7CritY8ENs5YD4Nd7QaCDGXlBwM3bpsrIegIIXDGUv+9gkI
GPLw3Q+AaUhb6a/hRJ6K9e43ZaqKHPHNybJMz3NFncJqJ6+vihRCzbm9ctWlo4p1qGW4X8sThflc
1qMjtcxEcPnXz8HQSUHZV59KTWNVZs/kmghc/dN0BKStS7TALmaAkKQeui++MVDOlK3CniiU4JSR
6vSi1+v5vTinnkeUvirkO6zwvPSShiyxpGArW0lgzb2PFT3rfb/g4XeBm04F4V2Fq+RFefq9Ps1n
HcaYUjBYJ0yyP7fKcEJ0CAjPjadyfbnHV6a8/Fi06AdId8F6RTo6nabV4lfapwJYwNHU3UQStgHH
/am6vvBmBmV0wusw7kM9aqicN2ABphCkihXnGihiVioXJH8wTY/RNkom0uWDxqfZ2mdXoReXyViK
F/ceEkSW0UYUjVFaHdXc0Dr8h/jev3TZ2mZnhANrZ3fksnVqxHurOE3DRxKDnSxTmSZkQ0USTSWl
bI27VQUHWDO6wFdipyE0XYZuHyAbUKxLOBuhZyL+kRQTOKHSfYJxNXT64yHW7NwD+ug55zw3ivFM
xEc9HbNfgeTT0U6AzHHFib+P8oh+3aMe9yYZ0EfMnWz+uLOKk3EN7O1ZZJQsDqT0bbvNHWKbKs/K
+xF5NgFfsKo88fj54Agdn+zYJjuy9HkOMaWhdRPilfC7+niDgNPbd3vH7G9x372ZbII8yxO9vk1p
6Tm4rUXUZaVfTw2eBF7hr3NdwZThhiD+1XOTuXIZeyD0PMJGNIN9VxuqVD+WEow/BuiO8Xmn7Yus
B4adXXIWr12HqNKQCieUsGl+FwVPPpih7HFy2oMVxoV5qVV3rzrOSczVCL1IfaIwtfZDGVsd+9Tg
uciigWYegml/Jv/bjUjq1ffXof+GxFAv9Wwg4Y7TDsOMZFkOdx/O4FybSMZ/w+zAIXLTaxDgJ0nw
Br+PTFi1HJLK4vhIw54p1sv+LznsZ1ExTeVpTC6fA5HjR1Drj95lO73z6VxrihKlT0tyyLh+SOfo
20jyooDgit2GekoUQgPKsyEh8Gz8DIc5D1o4yuePdwxKL3sehPZmqKU10kE95jGOaaYUsJq1/4Po
g9TLUl1Q7rar8vs7zoQ07yypVajoXtgS2D/bY6pMAWSZqXy3vyOopKu4HzqT0uxWhC7cPUaiwx0v
/JPv8t4eHexU57kVSrJ7m++l8EYXHXXZysZDvTHLiZNK48LKhIJOp12omEtWhQf8DOfI4Qv5bKk3
00CrJLh6mK3oGYzexagQDe5NhkVXhPb4AHxAbPk1dzfl+hhFr1hycz1SEfulMhslUXrj49iEyZWs
IC/rS6RdYh5Wz8DUXAL80Zy2zwHSuPpsH19f/U6Ifeb4EAWB38asULVv5+ytB2Il5sgVctcyvug/
Is44Muq6raMQfJzlYHtWSlmzuPVJUZeReDCgJubAjD0U8Na5VNcWNcykRm/m0zreIjwLvvlnHWtu
ubA8o9WIT7HCWHB+ka3GfQgSu5KPTZLm+XcgnRJaypY9vYhfJpxwqxIHlMNcMtFTG+mMoC8v/SRI
o13Jn/8OLr8V20XC8FB8QbEZ9OGj982LxDykXywmcurmAECJzzGgdiHN5Nyle1XR9wObZaM0mqbp
KYXTS2HU6sl6k9znL5FvnsipgocUBjmmVxIISZO5CDRb6AKbyKyFhG8JE46I6fKB9ye5SGZOX3Fj
cmUQAobp0K4xyPPB384tYkddkjnE5voGq2EeH8ftqY3R6AEypMKYqkNHH0NMw7SIF2bHkY/9dkzH
7fF7hJ2UsL0/7sk7R/3sG5zsnSWWCKY9RUcs02oMntIIcKg4gj5nDhYz/Df96Siapup3JDe4nRbJ
zKbuV14vMScrsgGXraK5g0k72ceWgc3hYv9vtNjqnEcqBcagKvVjslSBEqJiCJ3E9Z5047P5ZVNg
dpYj0d9Oo0VpHIjAlEsz3QEHiukjnc6I86CTjpcMyPSU9pKG8tWvWH2IFoYeg74cGeTFyk+FJ2ip
Q9LUq6mlj4J4kl9BBr7rWb7tGTfg/GSbWzopr1cnntxJKAxhkt1o55peTVWMImtSQkk41cxmAowL
TNsujU1mohxXQLFbQzhdx7Nsv+2eqadNZwvQvBSlDgsrkHScV8hR2dRaEX27wBW5G9hARuubGZjl
XiYjfj63oj4vTYaK11jP1QpyiSirCG7U7FXr+PoTtiWyu7IX3Of59klVhH0g0SeXYW4iQaQaDlyd
RT/127+U2xHlKCSz7Jrtd5BXF4YWiCtXuLqI1l+G3Gqqsd0cK5UvY+GCTC62INrxg+fNtS2cke+H
g8CNLwyTwc1jO+9UU2WyQHFIEwj2p+5nX7WdWl+Xp13kIICRRq+YzATYn6PqDAE+AqeIOc9YjIy9
9C7FfBFCz0Giqs8ms4Rnfuo/BtNWSqmTKXR0Xyoz3qnq48n5wdDTvbU90FaQ0Fb1GYJfRstLO2Br
OvDgM41P9+IBI8PKk7UWEwNYRPmMQNqKPyDbpxJ20TfLdK6yC5ZTJW/MtR/oRFDZuxw2xA0jmi7A
HzGG9HtFSZX0/hkPxMR/a8NSgZ4uQNwzf0na69+Ba0oGKO3kwUlA1IRWdAkryymKpFW1AScqO8gT
6uV2wsgGZTAhoMaU5IrWgZC7IdFAmSTQbfE5Pwwh2Iyo9dwqp2dOIyGDO/gi27rnkZGScgdggfSe
JgFqwQP1urAGb03bSQ8kzKcJwSkzWuXlByyj5ERDeaz/8URS9ZXPnPhC0n3BSsVXM+wskPWPgnb8
gLn0RHZ63YMPq7WjW+/+1qGkeKQFX4Vy9SCRgTf3Xf3UXPdR6N7lbtccKF5m86PE924ftGa0zZvw
DSwhNEd50tzT+9j0SYZimRq7Ufe69dXyz/DiSpfzg/zeswMxtE/feVdqB8SQq8loNo+ntB4xtJyX
1hOO8X1RqEe3IdJSwJJT/cIaCHuEwRjl6SluIOT2wRmb4/PGlVFFn183TuAhJ6WLrFBTlu1y4WfB
IUmz4qMpyIyHIs35VN1DFnIueS+kDa3oDw+0nHLaYEwhdW1lQ4BaID3mPQsvA/xsD8nqT1THcS0c
g9iiqPRturEzFQe6sMfh6lPsYG5dT4wxcxD4AX2rzkLR8NeJNLKVnred/GArgZXw15EJKufzwgyu
eBAclKBLwpwwLpMUbBie19J9iGIXgKH38Wfo+eVvjqYyZfd5xLHme1L3Q2JGQjFqw+dukDnCwfcI
5W2vK9aEsf/jEfYCppBGXUaJC1BebTEZROWilRvY7wxaZSOc+RLD3CC1dR5XLKijwzJFl87nSKN6
+dqMTDC5EuFq+xr4lKDRrSNfMC9AXpfb8jDBPX6QwQKeHwucFhdkltQIkyoE0Ozkf3pjo5BFhsbR
xj7VLCFBFSrDY2YevwOOfQDuI4/J+JdAXeER+CEeDWjFP+XZJ8TKM2ZbCCf3N0Q4nf4pmmRXgid+
/8/alo41/7OhGW1urPjdQ7Dbvf/KcM4BxsfpNlT7lJT96dvVANxw6viHkm4+ikCrzBPq5YcKviUJ
NeFVvCFcCXB+FxmPfwgaOoB7vo0Od5yd6ICf5vbrjdv1xZniu3UXD0nmBu50yvUH+IuyBBHptjec
SL8P9DjAvXvmb9Z04NE72BvIbhvwIvi/XvLG2H34zkJv/u1oxcqM2uxbkZ0pnPVa2wX5n9HZT/AM
sHbHR+JUvZgeaCmeNkmeZGCuPt6uLOeMgQJtoJ9h0Vh1wDASL57+ZahDbwTXUQrdBb1Z+qgdkxR7
gKAvwQMsLTR3DoflgcCtBozA53OcucjFTjJVkU/4iRIi1UXzEGAom91gRdJIb0jQNTp4fk+BsHwp
RHLqm8836iWJrPUJL1bbvAVERmDukmSVVSLzy9dQVq/GKMPBgXodwBuPLK4AyIFAX/YHLil3ECsb
iGG/RddgXuIsxp+kenAF0mBc1oHpof4ZlYN4aXtIcyTHwfQ8QrcbBEdc7M1OhIM0ngO6O8YGNLYD
qorwo+cxpK3LHuUKouQqY8P7nGkop64587RRP4RsslilTLOyFrDXhyBPKFpCp/Jfp6APvqNKNnG6
WApcLiMIvNVT0QmF0DfOxWzL2fEM7/fepH60MeexLgwVWOaTTMNvCIPvY4Rn0H/MPAzWnuqzg3/k
rPExJcqRiMO0wZEkUuO4yivAg0X7gzBlk5/oB9WguIBOC/JkzknYpBRNvA7YTBQYzrtswPpgGDs1
TuUTr3f8bPxKSHKsxNLDcq7WiO2CXVsDy/Z6F1g2EM1dE9AUmF6Vb2Lj/Nh7N6tLoHFN++cS36k9
+m3lR6XazBoQaEMpisRK+zihso5ZzNzti8RIdnp1YTstxfHRwqq36ceDnPR4GoOnK0Xo3Vh1Koc1
XVtjTy3VR/FEtacPGS9Fl9imzZ/paaVz211TU//LO0Z30MnKlguamTGaKZIg/mV8R20LqFYMOOsu
zo8QznHYbKmpeOLO9MRa4lzQC0oW4T1gOOnNNKJL+oBTrjOmLTUIlf3Q8YkjipGPWoBzSXWtmE2f
by6iW2tZlxqGDatw2x4O7jrC2MM36J29x27YcEWyLHITBuE/hg0148HExXVpD6wg6hCu7ix8gZOe
8BBVJDCfLblikmaoPN8ChRUrhylK8jo14Bbj5P+r86CCerMEwPCENFq5IGHvPi6EP0z73cpE5z7W
OIxpmuGK88mv0u6f9mmXSpzZj3Uxg9+rbC+SscTfwkBNr7gA4vimt3r3RXORZjekPY0oOzL8bmpu
i2Tpfz8VXduCnRzlWC+itZfeoGMud3yXcCGLvVFcXhfZ/qu2mThfb/vIY2qJSfJ6csLb7b9u7QxX
68mR4eKpgtzLBwXHOEbTmOgl77lA7Ey+T03wdwTa80oLonAAJ1/PmSwQ7D1d3GLAn+/0m63TuzM7
kbuC9p6U0c58cBTYIaTQ58P0hHeP39kWdFdQkPvu45sl4QZDEMLDhocrPfw9vEF6pqfvoJAinVkG
tg63mUGIQaBMwd6riomdOgagsjl0cX4dIYAXse9ZzC4JYQpjObS3AYWHAER22dCRpMfB4CXYjVtv
ScpWj3BXkjOeUITKvgFbcY0LnpoQkuN0UbUiJRP4USDCUS7IgY1odD+bLlE6EezOFd2qLsorOsYt
LbBPx0vVWEOfRNHRYDCOv58EXudqEC9MY6blkeAo7w06cfUSiyx3zXtuS2303hIqZ5dWLF1lersG
DftVFPDmKS8WaAeLa8AOvAHFGA/mEdMEt6Mt+wyizy9QnDuIjBd/l0d+pVAJtno8gH8Uo1v1rWz9
DMAJObMsRAdfsz5Fu6Up41kbZTlj7v7QvhBv3Dbbyi4G7tzvPdRMAdtDhb4ScysOHAwJSg6OvIBI
03f/olns+z6w0ca9+ZFSLE0MUHPZlaDZJuvANSjaW1g198i0JXxk62o1ReqXh96UkMxcbY5kVMZt
3qFCdvE4dJPYA3iT504NixMAnTA2s/HxG0rbrZ8jKJHWwiSB77QiuWxA37Nt437+6+FwSzyYzyEU
uLYMbxSJy3jVchCK9NznAEAiFkgv7gE/6yeIwNN2IPpu/1TV+nKZcV+zgkMkjlxkojjEtXDNvQhS
MFdplH2gGeBhyWZzetkn53AwEAX9FqDjYSzAx9U9xsgy+ooezYsQLdMzTFQbYPoOKPxztU2+FrwN
U5G0uS+r+JsOeXbwYgK34us5EPWTMk3qbTJMc8N2hLb324Jo8JRypfJkaZgospqRGybN3KvdiUhp
iM2TO0y8SWoB+aF8W8kNhy8RhM74yMnhmlZ6VUzfcMmtEo8utDMDonz0f1fS0EFJ7aDBTf33Oq/r
PeHeBRjgK7Ji7BcqSz1OWukXhzeP3DyN50jUUXUnzHUm4WVZ1QQqOUfTOvi+b/3OADbqQvSZAQMW
zKSJDUm4mqf06oTRtjJ28xffJFexNmPIzxRVewhhs+WDW7/rEltR8T34J6JVFGJ/aSrDNTx8lunK
84MkFwaZ/abGisJt089Oxv+ppUYRn5pkLGSOPGimqOyce8PwgzO4+ou0t2PtCPE1Lb8EP2ZxV9qS
xlsBYK81fQ70Dj9wHlk07Y3qPx/t8VlJLepFPVRxrFSOeZLgFTc6iWuNkD1p/xw77QSFANQ5EdxI
MMyKABNUIDOvT1Rnzjw9dWXd1MD51jX8AEW9nIXEe6SydXW1hV42dmdlchIIdAc+IaNmkX/ePJlr
1hZ6Ktp/dw5gdhuqJnlA0mzjEGeboGSJai90f2diG9aPiQLGXa3mdhET2EnnkUoz0BD9HSFqqigQ
+YdScsVo/5p4qw8nPlRuoq5pO5P3UlxFl9R+5mtogZ74laDrSXff2xiazo1Dkheoe+uPu6WbtgMI
Z0jllI6Jg//+H17Eq9UgRLtKCmHQU+oVPxXj5feRwwRzx6BE9IoW3nWosB51ubqt0XPy2Xur73FQ
t9+10D/49GKgv8ms4GUeFhfeWT9h7RLkey/VDClE6tJUi/uEbooulsDFV0kyZKChFSESSENpYjy2
MAjybvX84RMhyIx2YqXa7mzgPq/eEH8s7xBFamF067Sfuf3cIlMKgOBdHrH/mIYBj7pyHoZgygbT
xYMxRLxj7LFby8SxT/E+15lf8czllrVGz1TdOrpZ7NOEICPityc9WmaqZ+zKV3hOtoNotA/6BlrM
yFpzB3PBdqZA4eaYlCVoxBmBDcuxblwatkYxMIzxJ/Lm/c8TrhDpRyH9t7bBiK13ecDKJ+5z0KFA
J3jMJghv3n28yBT4jSckk8UzgIybgFDrae5wsfmFDxLn419BjqwlaeR9Yk61WZK7bTfGMNE5UAFA
A6DYzisloE7E+KcmFPV9fltVWxGenciTj8trvJoPN4nb9G8EjA3m1vz6AfPiH2DKo4oIemAEglrh
nPkJ92NV5VvAPGLAONUkeUM3+0lmqwU8Mq0A3aD/vHRyq+RoGOX4DW3qw4TWxkPsb477zpbH0O40
5CJEO7VfFz9ajKKGMEm+jyGEhLGpSDr+cWHYUfH3c4DpR9vI7FBKRvUCYVTKiA8JuKCKfPwOhbOu
jUAoB9H0r0XqSjj1GoNRbXCNP9XJur06iJrMkTqcYMcGO2bbwcfdYApKVjyeuZ02N6pd/9SNY6YV
rKxMtz7f/RYMPMY4nyPwn3x5hItr9hZg9/aR7hMiTk6yuuy4xQAsfmWdjS2rcpCorNsItLDOcUxC
aXMJKseSHTPERZpCrcsz/h4kOmyGbXB8kxnD8/WUETTN5U7cDmj7cFU5CNoPVWDcfAjeaKMNOYuU
ZE2Wtp4+UwF4ZxXAicWJLu2xMo75PAVUsdFaWCA4Bt3+LgFSFKv1zbtv6vRHxonTM2iGpU6jlFoq
zbD93aySRF+iUBsTjukhRo/kD21kiYLPVmn9XN84NcFioknxHHMxpH9IFuuyiRaR37SV032/lyyX
QcHG2UwrtfEtXeHhX2Qp71crhPCYkN1Qp0M4vzu5b/9OvTAHiHhxY7A6n8yg8lf7AsBLu5UJvpKM
5j5pAHbqht7tiohKgVbrm81NrsjdPYj98p8FsRENyIvitx3hCIM2CtHX3KYxgo2fttDLaHFEirn3
u4xjfFvMtturr2SUb65LWWNjDnXSwMarYjGZB73IpD9uetP34CU36yPCSFWQP0/hdjXEMIMdWHFI
sLw4zTetrh2bZS68cXkDpsqcNuwU8uChuo+rAuP9YpIX8P1amJ06mQmdczTJZwGy0Woa16Q1NgFl
vNRQ99qhJACPl39LCK/VFWf6a8s88XeV1zMFutfbP58xVTZYRl2DQva0gnvLtnxXFbBBxjFN2/69
GgTIPxZdED8yIHm8wcv6JrCe1GbJOH1BrZk3YuCqwbVwTNtmN5E3E59+eIAtnDaEWvr5RLimnlZd
I69/0JpIk9Gc4dKQcvGG2vdAIYjsUJuHt5Q3YH2/NQiyWE5HRD3izVvVOm3AtxNa6tQNxLH6cahf
GA+enfp/zHFZ+fvpph9nlSnQLUqJWX18US58PWP8v5fx392Fonpi0rE2AbkahrfHrWOJ9gFMJAl4
viHY7mB5/g8xOsIDV1wahyZmmCL8rdj4B7i2v2yECfl4BU7ggHNMKRXLl37s24GOy/FajBQHNl5k
9l6poA61clp/7Y+DzagD5COW1Xq958Stwi9NPwfBddWECdYF8vsucprGvuXn1TnrqLWotQmGTzlk
TuJAeMdEI9dje1w8FKKUbYlKS6Sl78LAq7viukMjlK6bQDiYFtuzggXV50BXD/d9vUCyu96I0kxU
iUbJQM8Vuyp+jSNn5F9UNSV0la2YULW4Q5CAjRY+e8t9NrDNMZDzZLS2tlr/j1V/EM5cJFrCdzDX
tkWxboY4xIfnVwnGgj+RjyfX+HFZErJQdJrQCnRGgjvCO6gk4+DOUgk3oDSkUda+5YDWrxdJz5x0
jAu7XJ150esHujfybl0FkpcauJOS07FTi7xnfOYLq3dBQnaPQ7tT6LwSPNpAZC+05SjK5XqlnslT
LA33GprWJULdoSjeN6xHvdzRNHCn1niFeFXgDvur8lxTZz98BhsR4maNjgwDN+2m0kxuBt/AcwJ5
9Mj1p6LyJmK+MYihWiquahmQv28p2myvT5A94A0K8zNDIh/cgtF3rtv6CRmVQ+6mgnfGmWc2Y0Zs
T9CY+qYwFblSrypPJQbA9ns/eezCHne6N5r0VelXrI1vsD8hzcmbs+NtxCyCoNGGsl+BR/we2kvv
r4Skh/wnjZwiuHmDuCTpc6E/iW4lVl7K447/OhG6yVF2oppdIWHRoMD5OLlEUFnX7TzeZSTANrzD
VBGhdIdPK5+DqzZ0wCN7YDpTjPdHaGcK8ygdFh6ErRwgUopgNbrM+cC14AmTBF6fcl+0aBGEyfaM
0swCsgsMkX+j55jtOZcHs0Un1rVmal/GaLaiv0UDIaDLG5wLjpOsgX9iMwcIMB04AuEgoa1hVfJB
ztlh8hlEmgkLBeQdg8VSLN3STCxFKy+3FKGBYKZsX0TV6yEv8AhfFNfzPaiz3leoBwvcN9tfXXzZ
N4czUmlrr2ho+gV3EXqnRB3atJpqOLQE5D0wVv9QSDG2WABsiC06Z9i4PGJ0teqVen1BATvBrAHp
TVdYHRbgI5OGmHjUr8Wbms/U7C1IgwJEfX6s3Vpc54KnwR+Q4ow5ksgkIxT8DfFYiiP/zO1LWlLD
JWiGWqXIUrmWDnfaVpBY12Pytl65QdGjxxvc463Rq9y6E3a6Tf6C0jXePbHsZMTEcCGpHSslZCW6
bLRgwgsNy7yU33dRcnK+Wk6mm31pIqZ7Aqpep5IC+KKOwHJES4zNuCDo0h4tRju1qZoj71gaEQ7N
f0tB1MdFzHs+ppB0D6FEldjC7+//pOW2UxKgsh/WKdDoMi23WI6UpkPRivrNsakdCBFRdEhAbIYV
oTJd6YdxYBGKoXo2qYSBNQ48/EMnvdz8UEKKBo9cG7Sic+9kvyiVGRHqWtK0ajEu+pb/s4xh94NX
K2gAFXEI3U2q0aOzqtz1WtOvdI2p0+vRr2vUMWU7dLymCpTAglIQBkkr0yil7bGl1belqsE88A2G
BZKTAcOvC4Fnn9AF4UzhvDYewAn85fVglR5KC8IOSL0sEfqkNG5L63KM4MYBrhLJ5KdWTAc1kapz
mySlhwudMW59h3a9zxyOapmLvB3y7FPOHfhelzyTWFPsPKLNf370VWNF96WfxtM8Vq6w4kusjUVB
OTc9CpGk658A/xW1U7t6r7QZd+NAYbBYyPMrW18b+BVZrlqifn/N05zI9B3YKIB43qc/1sZc5sMW
A8/S3XN82+NKQ+4wPxq62gmS0UcwS/sFzyG9qZuKYb0xbdzNYM6TbgnREDZk5vGGG8yRqmLy9y72
X13ldYYoZ0nOkJSYDUQnNLuZ+sU/hjEILaOI0UKU6N1lFyIaQYNdf7kBf9+4OPwJIZvOdV/DDdzH
4Q9lsgvA9C7CRwFB5y2A/etVkgnDh2muuE4K3oV0kFPL/qI7npGrmm8q4GMZ7KZLHuMJPITytbWy
XWyNsb02XsBZdHLqPld7/wTbDb2gFA9Yum0OGL5bxtU3noqL2rniSLHMfXarR4Sr23LdkNhRlPkc
dh3j+Y6tghH3vBULt1AJh5sMG+GPoNFF9WBrMQtkbSgoWN8H8Vjq0phZg24gZ2lyJYwxV5YomEAl
31PTbZ1o0j8XE1nugz8nPxLC93eTq9LCxs6dpXK7j9ImEe7CGhfDOyUjegMqoJn95DEpkcs4RYuX
B8lfslWhNfcuna2gkoE/Bq8HYQvcvFJjNf4Nxu2OovuayDwsO2n+RyundZHg9wodg/uJj9KQjnes
mfDrf32ejPwN2n3jpZMi20SOesRPRaW/Y5Y2pVCv50afSdZoAeBzWaToBlwJeOGNL1mnRsk98yl0
5eM6008grD80zA7OeqZw+58WKMKV7FJUcDqY8ePqY6nSseenoNGqUrlQF6iRTPm61mQy1C9AO9ue
9m2aJkgkIW+x9XyjuWj6sTlZ0MDYifZkMh3ZscwvL+xBKhqpMWQSEXzsNGfgMiWrhXzPaEfz+a8u
cKk5l2i/vR42AeRStEL7SrRSa4kUWj33/dcPYjkn+1LF3dgFnuWg/xhg85bf9olgh/xumX2DNA4/
L49wvtm5TUIBiw4tVHaha6mBie8XCDQ/QhCInQNgY0BY1vURB74/Rjr0qU8RC33ff0EziCZe4DXZ
0ji9qpV++hjX8O1fJAD/EhHmMhy4GVjKDEvPap0Q9Murf3NTRfa+CKbeIU1UGs2enezVgAOHMUGB
JXVn3YfcOgaaZRV9Jqg3Ec6Mq8JepsrVF8Bn/q1hysXTFuTfuN+PcloCI/0UAr6uSDFCG9p4zzWz
wPeg89/y/hpZ6MTUYukiPjmcGZ+cR52lglvigNNALd/pf3qxcBRgOoxN9nVQl6qBuggcKf1ZT2V6
DwN6M6QGHpXtyfMh+/BB8zIveAkeWLFxebX6K6oX2RfyK48BNuIZsaFT920WpOLik7BPp9Ae62lN
N2GXRvTNtPxdN5FVe4oW8eS3Lar/tc/5UiO8SqaLUoxudA0dsRc2FMzkP3Gatv6XpK57y4KT9QH2
jqvoP7Merh9vN/v36+PThby0LS7okqUbe44KcKgabhNbwtVSaZBjr5MpVxoTJnes3W7N1cEWkhIj
lvmCMD+JWaUNaR8hV915kR0LAK6OQeNz71GVfERWKTU9hryO73IjpCJuQYqOOvS8WVHfiqvTGAa9
51yyW+m5aMxKThSk6g2AtDs6G8Q2Xi5fflxHtAQZmiKhSip/rii7OwoaZRVuklQuxtLVoCwFXbnS
bISp6QltXpmy8hRy8YD8QmbfEXkw1y5J+3psWv06jGjo4NNVDWBs+vOKg8q/ggys3K80oogLY854
Xu1XySjQuDFgdaOvSSRmTzuKAHawf5MCxywhcchrq/XQOl9stNZ4zcRFvxpwHjWD+gVp6Itn1kn6
zpKemQQyp/dZHcOAUpoOn82sLd8/uuU5uLEXjz6IoU0v2J1jxdmhYJOkuz24osj3cdbzCTa6RGAg
2QkDOeT2wPxC0ktuxUoxjDyC6SLi9X0eVozyjkPVMKuV3rIpxzkRsGe+Q0ih3u7WhW3jtrzt4NQl
shsVa/kL8vunfIGs4cO/TJ2uL16Cbdc38DcappyzXJf3KsSQHOYkhvQkDjOl8eZhqQNWfsw58dxp
i4Gob9B5vWjNYt1bboMWGRmOagQ0SPIzcLGbx/qaWAYytBfjOAuqxwS65RjUryRLLZQrDKeiLoi6
HxpTii8vllEz89S55OZhfIFlz0VfkTM3KXmtWPUyeiCQGHqZqawZvSGIzs52JsVSVAXn1xoaXWNv
o712AUSZy3ptQL8UyWH9bl+F/XhrFx4PSwtsXKMGBCMSdYpe3SVHZL7EIuF31n+nXLs9nx3KQOlC
geS+68Q8aW5ciD3pXTr2Q+KHs6NspnTWDAM7gJDGOr9qmM/qHCFTfyzZUxHVJIIoqLp9eO3es1rx
QXNdQat7Yr+1q3xIfm7XwJje1ZQA3o473ZnwUpXC8clgCWUPiXmBBGG99mQ6hdgGk2DJ2y8+ap3Q
ydfkX+kx9VwzVKHj0YQLDlhBP2QGjX1GOyeCE/s0DGElXtQJ651TwgR47vOxiL8CeVziUTkDC4X5
a0mTRn6F70+4xf68rHSwnmScrytP1yuidXzKGH5MViBX1/kZpNG/XwAr0626H7Az8IlezasSF7m3
drHCPt/wIJjXctr5wVSVAM3zyBjasBwqHbMZj8/wLJh2Va2afeNE6CArHv6QTKGflg9KIB85zeKq
qz5mS9JDEGTZq6mboF2QHPH1aTfU3tk4kRTxXjzayvrNhuwFLnjJYELTs+r4AlGBYqbZ7KH90tHK
ypsv41H4igULAaFW14bPNqnujzf04ufylWa+5bHkacDfqoSLuSq0u0v5lqW0jK7uI7wr3T0pKPsL
lpdMu8z7LQfTUcxI8tGU9ROwkxAdVD+qUTxToYFpo10G8+LtQjn+kOqWP7Wt44e7z8+0bx4MOEH7
WH63df+dlxdWMLzKgNuoIFMzHrG7ah6jC3Y7Q9kKMy1T99yGv2veuKaVS4qY1xzi+NnwWgwhb94j
xR/VvZmN9h0NHIiOV37c5JhsLtGKEQEoGxW2Jf+o5EE0rQ/RVPDE7WebuRY7+Pdhzx5NwP918eJ8
eSYvBKzJKzDbSJdCIg8BDnsBXbpVHqgdFGtTsvKOeoKuL/2rVyI8JdNhqrdJlHvb6ALDMPZep3p+
WR1LdsypcM463m1F3CK0Mu3xyNiFUvRAy+xo258nX130IGaynhGN4No3jJMnuMt6YeyiTWuvYXZn
Pv8WObNekOAq3mnMJptO9Qb+UZKy7jZJRolPSoxEs3TiUrutP8SjMp+nGg0SEHYnOr5Yid+sL3ey
ShooZLSrFEC+CsclvDt4wBzGYdk4zJvvrBi2Dji3o1cIzJWBvi46BqQn8LuivC3nMW23zcFoNRb+
qf9ljuuQ3Z+UUaxGjlMSXeS4H1Ye42pA1fSfyAtYQjiq52zCOzaXxoqVPa/LFLB55IbcRjj32tDT
ZILRGYMFWf8uQws5Ftu0n/Nu9sv/quwqYbFFQoXcyWoNixQgFQsEhinJisp9mvBLAfpUD2qGMrx2
GCX3o/erp6kSbh2OrIK+xwhb6sETrXtwJb5A9qYK5bYve1jh6C5bSKN2ezEKVLNu9uQ0aV3HZmcT
VgnC+nq63tuIqo5E7ClW+Hlfe8gGoHDh0bLo7obyKRqiJsNjHyZp7i8hqfv+4fSWf36Jz961gkt+
T0IDGJYYA3h+xCcbzBiu6kerlj7bVHNGjsjRYL7VSnj4/dcgrB/iF3PPH3MUxzn3iHGdfzqKVBXX
kRLAkCnPC5h2fZQlQp7bCKLa0gaL3AsyIJ+y9H165bJSQMoEFrWU3tmrFTfjYIggemX8rOZMdsk0
bj/6x5Wt4M7BQ2mhbo7aLg9ycFgdFiRK5KXUrL6g64gheVnr3alkkRVC12VFlAj/tA4UNEIRUTop
Mi274FvfoqWDHqJ0RaYId6M9l5rI0PneBcV9UGQavj4VdEPwYAi7RYTCegQ5wW4cSvhFplwoI2xN
eJdAiUuekaB4evkStR2WPDKxrk3bJJkitiPA/fp2JcVWPZxcJLb3sIpAdJKglOrI3qF9Z+C/9b+w
VWw8YgCoa6y5Jt1+JtfpQIomc0v7HM+lYL1dg5VyKTK5p8IO8tUX5uNNZ8B5wGrXD3tg3K9L9vJA
rOfvGT2YE5RJLyE+s3x5cyS8rS9Xoc8/whhI6aOJr8EGPIOEA3LKW2GGPiuUnPFh22WLUU46DQQq
McdYuord3+XCBCdLH8asO8hBTgIwJuYH0S95IYTlmOp0zyt8I8qtEZm6f81yL1vcLkVE/q4xHKM3
HHRUjhY/bu25pPYPOGnqtrnWe+pklJbbeLXcpF+D+fUVOdN350eJpFWS+fgk/KXuaITjgZ3+TnOi
EBfkNIfwEqYBOew1roL8Min/ctc79pW467BnZpvbqHdP1x7BuFx6WuBs5CB18TR4eKBsPcYS2+ih
GY4psCTf69yll3RbqxhUNNO3gQr7A025u0l51PamHvU9iqhfaICb7/Pg0WmO7C0XiGKqkq8Q1CnB
R7qegzyakN+4SrcDJebPwhih+ZpCyaGWcV9T1LCO+J2WxFziGLL8TpyLS+Pp65U6sYde8WAKMzS8
pfSiO+eRdesorwWJOWAIcvVpJGpyyViTg1+BCpbSGxxGh5a9MHHXPuI4AvFkeAKvmEgBhAnvlc6N
GCsciZKND+wfUlpo5w6oUTWdtH8ySHzjeAFDNDfTT5tdh7BxdoeeJHdYCF/BjQoWrBY4LIOcjesc
4q7F7nkSw+d6ZHMYdYgOk2xFrDYGvED3bCnSIC9hU/4PTv7QWgZaq7ivf3qNlChC1tgXsL7ZLUp2
e4VLLuAnUiTy2ZRhF0r+duwS8tt4YVemqFRK5y+VI/tbsu3iuu0qKYRoA8gHDjhzDBGVZSITzp2C
7uySzWFxvsKPhiRq7v6fgZ6Yj5lLk4KXCfrkNAHh9LzmPKUgM+vz2GMFwVwS26javb3w3+I+l41w
SNNvvjzH/B2kt0A/2RkxW9ksO/XBK/OaZ2lDUqIDR2xgPLGFoxPMk+HXzgMBXanh24upd+XZVDGN
l9fEDni2Jf0sB8yi7jLCAJ4z/uDBX8dmT5/W3BTfrgyRytzSMTPMCO94nyUzCDWS/qYhJx5uH1lH
iXv+UzwNKxrlrh3BdgyAobGCSWcFQAV7e/Tia9UIlMg6Xjv/6ZGgya6SP3QX7SwWNuXTVYpo5jg/
KYsgTAlUVNGY3TO2vShqgu+tiHUYwlaWqtpaYvBU0WrQRszUGOooUv4PmwhrYKCRP9MV0v7dQvtt
lW/kCUrE+u7x0AG2yj1EIFkmYKoTtWir6VaTQgvnfZ9lTV8jvwysFTrcixD0v9+TPhmk1nRKBg82
Ax8fYO+AbNK+Y9xmi9e6oiWqrFNCjKfKagFDZw9WxCisT0cuyaI8mPxYuKGW3XQ9godobfiDcqbu
gwx9xPTvkr1BBlTgep1ZOuTcMi94DXz0cyP4m5G0Kbcv4UdqFmQAZ1NBr6Pqq9+JXML32iIMN0+1
d0owW3ZQL98yODkcMiR0N/pz7HTc4CURjGUV5D1nZPlv4F+mdI9rBJ0EFzN9heWBg7jn2yjC3IET
EdwaYYfrPWFq6pdrxmuppPBbx3qsirCooWIB0noexYhvMlRvySdfppCzxveY0Ds00ERJj+sHvKrZ
xzMaaQmGJhDfCW+HpxigIXwDdhfq7TJuL9M1YkMMQAze7Cjfn6cnae+qn6LKdv+MaWx6Q3NnqygF
1rdHtBj5aLggfiSJi97JNa+2RGsM4bGfeANXDwO65Iz6M1pLqH0q6U2mNIFHFZu+e39xPhTiBxUM
7xb7M68NLr6B99/lZNIdKM/G3wXDPnTOLPC/VXzq6jPsHKV/bzEJDwXzGwilH40oG/jObgFj1v1I
UJR7DdMge5m+M37oSyL8vKF8YcT5p9WfjRH3SS79I2m4WIh0neX0IvNza+TNzVDb1ko6hHovpTXH
JQO5YeuJllPkskexc1/PA1bSQn5yK3gtnflFlW0DYp1G0xBoThevrL7nyl8c+TT9jK/DTiHS6kx8
uD5iAiG+83Qc24DzPSnYnE49lEUM1VEwt0NEYVHK8kNfm56BkNl+ZvQ6DD21uzuvWv665sPSzmKi
/ABXJZaJdhiybBKK+sZ/ZyO0385jy/bwiZZEbSTfqnhgd+Xq9OlyBOujtzQhoylmD3C/JW9/CITt
yMryD6eLwTiIrLxF16tNknAyK1EuT3ui5SJ3SYdEMl8/4Pn4t3N6BsP0XE/o8/tA5GX9Xc+Jl+Tx
pbXhbSgf14hmjJQ4GidVuVDBTn12s4Sl1lw6MS4hbZzZVd08ugaA72ee+c+98cfzl8oPJyRy2Bqw
CnrbFpl5rNuMFQ05cMCnn9ATGT0s7LUYWo18O3atqifkD0tbLsjmTzwyr2i57ka27a3Zu7GObeOR
ko1GW2jlGdDkmdpqrYN4EYiB5EK5CF5OAPZkctwqBjfhlr3uGIyPbhDaQ7PsJkWO5OJkYddrxUpl
w1Bt5Te40h7S0dhFbXvp3LEkfCvwIaSMMTzWpgvNDgyF+YqHW5ZTSvO/LXSkADd6nU4S0L+R6epr
i8PSboV/QvPvd1r0Z4uhClNH+BKqdtrQDQ++drMtUdNA2iEbj2bdx37aDQoMQv5yph2rxkAKT6KZ
35N/6atVtvUKMcqMsPB2QjHfFmuH54FXqIABLePktMYOfB1VhysD+ZAUP9Dv5bewnNbhy8LXe3Xe
/lLcHV37NkO2uEdKpn/GwP6jkj8uA5hKMYff4tlJul/R1hqZ3zVZPZ+N0cMbkeSVXgqtj0FU8b16
lYrJ5P0QSGrpk3MqRsFCzIyidfRfm8dkOA6fGB88Iit01kIoFYzqsTZz//vADVr5JdK2XL/+OwDQ
z6dUfpuYu++FpKl4I00OkuS91Z18dMhHhmT7eMCqCObeiKfylNUi41WZT/D0ZPjUWgHpqQdrd67t
IWtTnf40DKCWuxn6DJLioxO5AduXI81Dmhbvs+fjy63r+Jhv2h9pfsIZyMSueq4Ugd28/uvO3wug
daDHib/2TbxIlb+M+hKakWRJ2qiNSA8QM/zfr7dSjiqoHJmzcVwfd+vQeOX0SVLiopD9hOhJPsGD
yemWGv0dMG9fE0hmrEgj6I6F5iUwm5pjnvcu0gTBRk6qzq5++5+D0ffiQICVklkPiO47/5/8ut3d
Xal2C4TMZM2Jrl3eiCsv4h22Bmi4z/6++NZGeePqlbPdr+pCMSnph85KX5FG6YoT/yFvvm+ZVgdX
8BKwoYB3flJErnsWOkLn+njanOmg1B9yko19/oCIrfdlttkhI/BrOd2pU+DUYMbsOa4vazx5T/me
NHLVZNpVTSfEARYIjbl6mjcOn/RYieiP4vQYyC5y97z9JrMIRQjv3KYRz7fbFNNm+ErqxOFZeBcZ
8nVlpz19KrmB4cTUA8vTF3oBROHGJSO+6R4tkWzwS6oUeQW4sxl/4mAUBgs/tZnfFI1HvwULKzTg
mR2PZaeG4xlr0zrjj0496r52q/hl4NVlpuB3hBpPw97rGDQ7o2Wjvlu6sAyaODuhZ2y1AzayEx7m
YzRKZ4vMJrYp8+2ZYyzapKU1lX/9iFcxbS1bYF3rO2oXmBW7RgsfjQWXsP+M+dVAK4OMMNhYosVU
uzWl0CsfBEDANjTzOPGlvGT+a0Z+RPRd3UplD4ObdOhm3L4JVK87bMIGFrVTrN/sRzhhs8oFNY3Q
Wtg7ePazKThaeVWxlPBXX0Rv/AgegqmNoy044vVVpnYhuhPz2+y/Ss62tfqLrMrXN0W8ddpbEWO+
GQcRxSbQr8RGCntd8OgDIbEuBvBHJtyySgOyK9QtWMJiUCn1pTX1DK9d95BeNzkoSK1eOASFkZdY
eq4awViOpCnj3pa1y9Hi+PEdSroafxREeXgkLkoxOH57iWeEiudSbsbPukl2KqPL8Cgibe9bVuyj
UZXZ29jw4NiO934av3O4Mn4yyWRUQcqJ6uGttvNziSEJyPj8Kn1j7ibx9+CR1AJ9TGgbnFZDR2Ed
QjOT4BXRKOT5DBNk8Kng/eYz+EvcndtkdxasFQ65aUy8dY3j7oMNrMiqyeg37WJMePe4ReCzWa9p
eiU+UGXB7HlmNRF4Ck5//oMubbXAbqweSOhj8P8MKjVxJhG03jYZ9wtUnizMjBhZEVTzOWEQlHIv
dLCQpRzQVFHD7MBbVnsQYcn2eCYa93EjzlhHrdnoza1WaxgJd2GP0e2taDYPTnslMPj+dx3K2iOv
P9E/hi/J9HqAvHZ+lDl3oO4tpkRWD0xay9lSxHdcjsA5RV6+3wLKfnd7nPIm+m24i5ToY6MON+By
gtizpTT7jG8pLIX+X8DThuV9OmsKNLPqLTT7VBahm9KKZjnWAAHignUOjoZydty0EIp9alg+Q1nh
RIlbm+KWPirdcI3mrGgEC/F3fsvQNArd4TNOES0Ecmc2kB9t4iXTT37zM9jQVrulhENP+00eDmb5
5Ulc/lad770ty2cW2y9csHqkOjyF9Nhj0wlhUVyzftJSMwpJPBKvSSQGaeEp93bWn5kdAbchv+II
tpodh6e6votMXUpAbHp1pVSV30TKeRwJj940F6Pn/pUzrZPqNSyve5swqQVj8Fai3aYp19vqGPc2
1LUPQzpC084ocEXeJl/rmbUPfokxbu48Ixpbk0RumKsfL0Q6RILXxoTd1SVYrLeryjpHpQZqPNH0
WE7iqitAagCd5VM7GVKnvcNBi2kRBSHVlhgOrmhGgokxr2wZYoLrY0Ai6mbFnHeibc6UXjaTGxoe
0Ymaabx855WMBA/rP4IxWWZRs7vY7wIx5vvGnoSKPQko5wNmjSmn73sZvNWgXZokK9LkB2tAIpfP
ntpCk2G+hyjp3TQqnza1gWB1jJN3k86BjRL5MqXpSr78cnIrqq7A0vuFZq8K17yeC9D2vaI6Hwl3
tVr3iV7sUqNz96g0xN6WBhQ1BAtqbezLKM05Du8ZB5ilnFjTIevYSOtw7mW6zlEOHKS+Ap8+3/Hh
A/jz3EdRgEb7XVVrkrQuYsECErtSzQ8RaM7zC8sxBX318rxZxr0KuiI/2GgnRC7kEk1qgSCYOro/
gambEQMaddL2qAiksatNPrGYRFu0asl59h+eIbEL3CtTh8E6Cctyut/MBKjO6yZg+/hrVBsoUthr
LROBh0Vh7AvZeXUk5E13zZoaX47nA8AaEnBIIJlo/qjxBUJaAx7mZOvfhGLHMijjsSr4lLwitTKL
Jkq9sg2TT9G5126EGTfc4qQrwyHO6S9M7YywQMPaRu7Aw3Gx4uR8DRVMV8hq1rmuIMjzEg//nuuj
SUoQT7XMe73vt4mXC4KAWAUBBEgSUCTLy2YsOCGq3/XmndxrgvPBedQLenkyLU2T8UJoRn4CtjiL
DeiUO7Rx8a2pQYWgSOB3IENChWGIjB+j5x2ZskaE78pB9O5QAueejt35D506hWvt5gZZ1mjqrqQD
G4Y7Ij1GTqsdqFQQRbAOBLTxgXvl6Pj12+NmKNptwmWRHXALFXlUE3JY1nHcXX2sk3kwvDC0osWP
VPXLDU/6y1lc3PCU31oXSaPG17p8ll/yu7QDgWbscHHm/irIpDiygZhE8t2GweCNRyVEks6QgikY
qBgnWWphkAzaq/XdK9UTeyQMb7nPUP+Mjvr28F5QQEQHOkAKzmRRUypGBVFqz6MGrGh55HA+oh7a
SzMLGAPjf96X4T0H5Jc3CVO2aDANj7DNUlCYneCPEuB+O+vooFomDs7OjMVEqMkq2r/UHppuiHx3
o4T6Qggt0zCVHK7xNX42tjmJgiwDzVjV0XWvI6Xxh23+Vb7JFxiFEPMFq2+ODdNlY8pgRIobhdmX
/99T/QUmQnBf4bl8QUwgf9ss/qDdpJ0vUDk4EGgULOGWKySVQJ7dMtKEtYff+96uhKC8+qnmI4p9
ecMCXJc0nSkHZxRvMejq9KsscjbEip1kxD2tJs8pLKrUpfZnlV+1O0Ddkp0BHSTOtng1zddYHVx1
7a/jV1oZhoyoY+PHe0qUe48TfE5G7zjlwqjg0mSo6sT4VDTbfvDppubNgkvsnzN4ffADc/fkQGlG
QMA+tOb+gTlU5WZOZbF06xQg45EmEzTqIcPdugFAssphHMUtZ5AcjlORjYyJGXzarS+lz6QLSRMj
eUEhcrFRc5/dgz4toqfS9uTQhQJVWDa3jD4UkrBdo58CirKyCBZczC2wJZhx12oPKdF+ddKg+7KB
7bUKBTFr/GGQ0zBfklP+chy1RbtG1M9iqP60YDZkh/iOJjHpAX2vio6vsa92Nx/QgPZbKJaUOHZT
mUv38uMf5BFJpGVDQccmW1lkqZlXACKAThCIr0hqHbz5Qmz3sesXmyQiCGijPu9KkHSrIRHEN55F
zSAkHKOygh9ifYkKqwUNYESx+uVY3P07MSYxCZYjl3ccisO4RBOw/qiBEAomS2CeHrSMWXfh2ul2
W3etCv2k3rMf1AWNrPcAZD6T6nfXVaLbEnMUfUOoIW25Nnkn4iYLyQJzkRzBOn8777Q7i+XG9nbw
N910M6P0oXaajTuLi1Bj/SmZ9Hn8oq27N+5GylZClSCt6nw+8ABHpPSdJWUcqzvEPnLVEB3eD5bn
Sx0BDm+59rfzWtEAhRXd0S6LaAmuevLS5k9zc7/9k8ADk723e/LjbjR05d5626R81c3SvziPFOhx
SrstHEB/tTuhPojncLAYoCcn74tXXCoUMAF/5bfUl8Hzt44DaMd8gpyX9aPuhoi2Dt8M71FWbxub
F/lJT9auNYD3obDOh0MR6al35bdLH4hPS1ximAPAJGtnwjyahkxFXk+LEfJTDCmVm03Rsa542Y4g
/Wt67NB8Q/xW+qr6M7kjINQox5sizE4ikcgHRHy7zm0ZNBTYNTCoDv3hKO6aLnAfjq53bjF+rcNw
rW45PzD8pfH7TPjW0uGz4w+vmf6YFkrDkakCr3Mh4LZ5GEVmqSb4HdDvQEEjC6dmiIinmqYGANpq
csxjaKMaBXSal3UTWGOozf5pwk0bBqNraEFFm0TUF3fLK2+t0IIxepMUCM3zLe3Qq3jVHCtM1OE8
pQOpVqAxAYiB3Wv30Dae0zD8d4NiVKDbgqJgle3wRzSATqCgMaeOQ0fbLQy9JL+JI61B0XTJ5tIS
GSa25o++hd0UwUg/7w97Y/0iJ7W3ryJkLtk/1w5mcXoklvOvJU1p7NGqOPHKpyQCxKvXFKITb4OO
3757AaCPZol6rBBIEMyQdOtmZNXERS2BUWBAR/Kwt9P5pNbV0ECFKMNruFwb4MwZ76v1UGsqIELo
xCoWB36vUfRv0om7Y1orTRBNqiVf0ea1uKEKSoulmlwLcBHCYWDJ8B+ntHkYZsA16oURem2HyGMf
YoNisfA9C/YkkQMJbSge/u8TsN44W1kPXMsltkE9MkJyjmV9adLvkhUHyLEiHsJ85TJbxnBgn0x+
dzD/hLgkJB9q3lo15omj3CPL0BSeJu4Ny8SYZyVRIg0bASe9zymBYp8Zi3AxmW4El/yJfnHcNjEx
mmIAlbKR0R9kFWqbI+dDYkcOt6hHO3RV99z3g3biCmsaB5tFPaDXhYRfqH8tAN35BjdbySJxVwSN
SOYJNWMfCZ3K4rOgQ3oyr1g5gnezc+3qAB0WX9kvol9YBeWha6sxTg/TE6EskvM1MjE3O4SO04aQ
ORaipQymTvG9dAYtE5FHMVCp6HON+hMNxjyQ5mdrzVUJyDLuA3TCmlqd1odAOnAD9aFAR3McxOrT
XlA5jNKjiNcbfZNoWrwP5dKL50Kyu1ARVeEQAqltbVf/OrjNxREFwiqR9WYS4Z4ma1Gxn/CItw6t
Y5WOk0lTK2vdGU0zbzj3KFhrf5TUXiGRN48W/wJj0KQwze+ns+/TaA/N8jXkEGd1wwDjQDa1IYmA
aquT3mqpQyBAR4uVSQ9tcPDeUpoppzaIGX+XtSSLDDEStNCkV6zv3yDeSEDT4stqUcmvRZ54A2dc
q7Y48jbaCa8Ml1xCsDo84HRMZu4HVsioovVAgbuW+PsMg7cvdDcPrzKoi7u844HlNUVPbzAgQYF8
/7FHsRr4mJdrx3ZpGK9ohWSnhUXzCOeOJUPA0TePLq0SiF9vKYJLfrWuo7pcCeM9IWKqOV2nyGex
6w697nd8sL7gpawLa2Tlgz1pFFPFDQG4nBtzAuGBXNYHnjnSiV/7sIEYMmSt0remF/NvsBv7R8dj
oZBehhG/b+cfYbODaJn1bdzNJInMo6QOqwwtiGSZDHNwp4kN64hyayVWMjQF0HH/0iYy2OBm0JoI
LLgwXitGXzX2Fd7FgOuGr2dmUpKFNpfE1gJBfkGr9SdJ9mkfyYeEWKB7oGmIn3FVHl5rhmppSFsY
UfVUfRioZcz0uSStsxMk4m+Y35VCBHNaXx22SAtuzbFqi4mMasuPDvB1HwE7JGJvanpNjSRJSl74
JoDh+ckx7HSvyQefawJrRIPekawzFpRxZf20fL7G29BN05i85gAJnXzzoC19QBGkrluGRxIlIMrr
rbbK1KpNUtXXV/Aja0fYVVRtvGxNvwChAyspjqhAOMHfb4U05u+zNbb4weeGgrLMnroiMPhpVaCe
X7z9HkJY+8PkxTu/C4X98fetMIiIbVrtWi/SovEwYH6xZ9kwC8w06LKpmpVJ2VAIP8WqEHi5UMwT
DxDyZsLdu7xCwL05HeLt4np2r4q5rAYKkgXlaKNF7pMxDaWaVLhh4GI1PIre+W87pHEJzN42yF6O
c+RTmiqnAkRdSUQwpToo9bMoU54jn5FjRJhNwl85Lk6gk5bQWYBhgOFeO/b8/zUOIGnTgpSwwcef
LBgV76D5F5ZvXaVzV79UmWhnoO+r9XVDAAuub3U15VuzzEYQJ+Rb4zYDsXk3lLwnxL3qgQr9N2lQ
t6RL22C3jsZ4iXm4MqY7+1YQ/sML9xbZ5ojfG2o2nnccwY/8PDf7kW/5Kk7h4eZsKvjkR28kEzSp
vsBZJVa6RA+jHzv5yaWpAswcSu356ojmk76gUfBAta+/R9XmQyQ10yJGIDbwLRHy8D+aQua7rHP3
PSWG3XxNCc1ZucONukATTBSjt2s4+P8+y90JLrX+dmD5gP8TgB+FFe7iW/rBHTJEmu5ZDWrRm7ZB
NA0F/7jC20QBAqrSyuSvTRbzbOcUXkxF18oVQ+Jy4cCxrEDZBgzMQ7ZVvsF5xg+LZRK7hH9vXj/r
CbGfWupw3rIcbmHgriF7qv0V35tIm0bNkS15NBi4RXEsTLeZfxCMXazxmLDGPja2rAPjPeQ1fmxS
6GzYeyvjSgR6YJ0SQyBSY8QIHteC5dY/v9aF8IZ3uxRXjjlRNTtmlQJHlb0l/YokWZ5e5hZZG6g7
n4HjmpjS411B3DTobRzUksMxZSfMzeuxgeVTLH+JTTIRhXYJDJWhwpzr33TWK4XKPw8MHJD0Q3Gr
ho0lSsAgxtSOUZQm9DGGS2+0r13hsaSB3/vg99QHz0tXnAl0qJ4dt0IISvp0zFSNU7TKGttT3HiH
YPusMGRySZFHEfaJFUYILrfvg5NdOu8myJgcmPw2zU9m6f5LEqQ+Ku6TO0jX+OrPz/F7b9AQ6QwO
c303t0zqVVByxtgnFbQMvVbpK2b1S5OwgQ0RuC4qXUEbCP8UMA8mSDv83lQ4drLQqrpo1eNO8DkN
w+KKKX1QcBNe/3MEEA3wwx96f6QzrZk6OP/TGa7t55M1ZOzpMOC/DgUEex+nOsor58ghATAJiua+
6KEIBEgRzcHU4eoR+bTLChCUUXDKH5I9g+tCtHmmaMd2uO8rjEufTm/gYY2YCtVrDuUyfmpDjdGP
fQus0IZg3qwkxZdq03Ce7ZqVC9lePLBRKlAVGHtuYd66tcT+RLoCTDhEVHTN4oxynaccFetNckd/
+azhoefQVVJHfvp2IUL5rgox2YJzz/6s//DOBD92zDhJE9fLnGNnjjs1fpKe9ngRif8hNQYRY8An
4to7NIj+H5KbCIPjgfYyFVqw2EqGhJ8jv2kFn9p8E2JGyQx1/y/4LxSgdYMargJGQoAQa8I8ZYg0
zzGzfBpvdiR5LSMW5LOPGZ654cEIwhJqHxzrhivHG5PSE8Ppt4Gs8PFcfDnyMWSIlztKgLcunIZ5
GJhEf3NkHJ1S2zJ4b09DoPiRHyU4V0cij8izK+NeLrCc/3Nlumywxgl+Ky1IavqzzXiOxtnrNsej
BUBCT6WMQnDpJMKCRVZl0JD6iRMVcEpGU9Nog5GznCMY5j3fOvy2XkFeKaXvn+w2KIJPxRaiDQGp
5BFUZFpMGN42rWZTABV6Yh4TQxk8jREFErPES4EUt7z1a+xZCh7FyddHZgrJLk0WHtJ85p22ovNL
+huD7tsfy7lYnSIkWbSU4JFb/cOwnu4noyufgrq/MlwI0PWh6gt5TSiTyDimletY0DOi+/JET6Vr
vanCp8Q5B7zOin8H41pppBtQHt51KgMxze2wpfVzwBMJwfWowDSZgrStEmGC3g85AaxF5wBCCc80
NKoZBXh3VzAd5t9qp1R7qjCIWJ3E9lWr8HWq3oxJuzcVQaP2byzy47ilAHuuyxZp5ftrwx5tFWgl
aScTa51gJmwYq6PmrtZW11+znKZtda1J6B/HHtKE6flecpUpvaDu3U8ytk3a5eOk0vbx9EB5P2nV
qOrQhpiL++D2G8B3FpMsaJCjzOLv/o2TisnTqgvEHqmBjoQBSr8s+hXFnu02CTsUs3P0hn1r6GzM
l0dOEf/1DKFcWiZYV6m9VkhhZNv02kdfez/zMTAfAxzI1wIs0M0pop8MkRM0qna7npMHhmfaVmqr
4ZlJGgScVjF49cdJbtCdqu6o6/jlDraY9JQWjSG/yUmmo7aKI2OmYX24DL5yKgsDLlZXKRv+eBnK
qVRDHXNpVDqwTmbvzYlhIxQ7lsA4vdOEAEMXIk/dWUsJ07TGgJoLJK3PFpbHmF2GOLh9GbRM1UUf
uaYr6Nhcz0euyh3YQFFGc97veE9O/uqsLaj5bkN3QSGv4q6RNGQ8niCAhxpKSKgFXymtbbzIL4nZ
clBBQqf6HaB79IzMX5ImM3jbHbfEeOZiS/t3vtzV/2z53onrvNvC5Mt8TXqrkrrjTC6tMLwNyEpC
x9A51eLjUS1SzuWI5/axTbL2we8eBNX4R0v2/jZWZCIyaYDUPAoJ5Vu1Cp5DK8jKy306qpuW7/4o
aOjPUWTMB/cjH0IeLxj7+YUuhjkgYog2zW7XukxgJ2k0wK7AdFRbNV2TpK04fNRS0OaezHJbK786
cXqEmdwq2oga2GawyjIsQQ8awQP65BfqjCClaNSBGiubhf6AUblTqE7O5SGTZ5SkS9Psyblzh5dc
rz8qo8j397T7BL3pUWGgZdfDByI2zW4fMrMLd9lkWlrUwnnduLgl3I12hbmmiyGWwRDJjUiQeldJ
OAYtdfDrUgjLFwrrsfzYluzGo+08V+oFfHn62ovaOg2/epQ7RG5PBHkpUODZ9tUEcnEMrVL7A4dT
x3Pvry3csN0YDx0EDyZQhzB01gXpO5JWkCxzTzVmBHM4hij21zpgEq8iN4iiz7Hn9P5n7WkintEJ
8BHW2uCQnw8CRrU0nRM9WmvnUmrRX+wPeXdCY/c09gUmMGJlVsZTge16W1T5fFDUUpCfGrgYIvpZ
R10cLfP5UZ60bft5cmPpELZe2fKFb/pwVREVjzVbDusAULjTRlQYkh1NDtN0KhoqsjGfyt8LG4qV
oNnOSH5Fz+a4rwQF1rNRYIhve2yaZcZ3rHsNNYVCrHemdKtD4wpGfWtsY8jSo+IDW54HdWG/+Kw8
LHApMGCkzWqur5PoZPcdxnPFf8uquluL1odo/oUUqoszzWdKMPaXGjQqJdXSmJd10l0za3SwugL3
27TRHIK+7Gk2KJppt0F91q8Nj61UZ7vJkmztQ6tVOPpLnLFQGIi/vDu75iD1fC5AeQK59R+uVFyr
A5IlAQQ6yYgAEGNqSmLOoxz8f2OKwJHrEx2BZBpr4PDehz25EHQEa+g3YZlBX2G1ZfKXjrbzhUgd
S9gBLmRW+jS+ahRFR8IU0RHVygfLBZ6io26fR996SRiMUQly9oF83RXPCjC6RD+6lwgsW+8Kxu65
t8FaIecWK7j6+2w5ihpVCwvIjQsG3Fu//CqVZi79CSpM+mgrMZXK8uGJE3vHDVHEn+uAVL4oj96V
v3r3/yBqLsb4t35XHIlc+N1JjVlmprS5NG7uRNkytJ9cJ+qdlsOcvSeM9mbRxjwk/3pEtJfyEFVQ
TjQNfUQXj2KXn2eo+ASTxhImWSKVVuw83JM1cWyTS6tKlzST2wbM8B/OWkj9Sbgqw1afNN2Ky3I9
iCHNww7y0bv8EyITULzdtT6hiVwXeSzrCko++hadyTKOLK4iiqdZzUzDg8rLwYiEzGh80aKd3Crg
Kbcj/cyyGTp2TGp8KipPnhAYxiKp+0ixvywcO0P5JdofeK8QgbaZlRa4Nin+1usoLCzjz7PEO/vq
YyEo/+ApfWgMfwHoHxpWyRg6INU3GekfPOWOX+Gb1luvKcqRkQILKQ89J2eloA5b9xOVBHxZMS/E
GYjZ8drI+CHCSfLtJBYmqQXqiDKg0Kulr9uu3h1R0EIYal4mY9ypJYZn9cm80b5kUWffgbdg++04
Zqh5ybfvrgd/Qyc+L9YSlgVIhwB0NZ1x5Rhbpl5kSpBWbWmqAaA3HsmAuLcm/0vRaGJ7PW+ueOH+
C4GSapU2BqwTZ4WBE4UN2hnMQTpsUJhcM5zg/Jq3sbrA3oGoe/RlAKD9NOjtcVxlWIKOmrjLAk8u
403VHLU/Uzoa9bLVfOioO34lMdnoYHsXXWcVfpShfxncFFr0jjr5aQQRCOiEceohXvTSqqhx1PJ9
EXJX8Kfl8tGjkhWC7v8TY/jg875zJ+gCwpT7uhIXweGKe68FE5jJvePB/BBLieAC7UmmsdS7cAOy
KEojZk9TgiHuGFRp80p3tqgq8o3QXjDkJgXQeM8ojeGWz2sOfwLDn0dDaQxXrSP3KfZIBoJUAl5f
r2oFWS/Y4oUukoCha1gI1sUv7yNIh/ctQgRiwoW4DhuDn+3c9cDMF7Z8kBber0XYzhyB1TD02ltB
OCuYOVnFE4dyqTt/zFc5A2JnSfp/lJi8fYiZC5LV21ttI6ZkDzIa6j8Fxml00wUdpeuQ7SgsjtdO
UQyjTVEvkQkE1cY6kpDePKwHgTg8PuxYqQmLaA1bB+fXjLTAOOJGFq31Xyg88aM0QrT/ic6lnrAu
yv2FrBlAQhFFX1f3nACVF6949N7vYUt99PNR8x9A5dLLWecak2N9ww4G7Nx47ueGinGUijLonIBp
qL5lwPSUuOFUBL4jgJj5CCM6mWuAqGOiVWMI8dyJCuDSWBLp/il3rIeKvkOMeQtGGjkQyfjIVi5Z
61gO9sLhbi1ITSkxjBj5ceF/a1KKuuckw4Yr49mwbwsOdpywx0EQn0XQajEfB6hXad9MSh7zZ9xZ
8VLhD8kjDpdKCB5xhS4Rrar4Tbt7Sgy0sO39UO6uQ883XEDt3kKsHiSnXGw92Ndwo1o1tvrfL+S2
B5W7x/vrbG512hnnzS6VfMznHieTpeoYxGiDe1hCcMoU2JSQHeGd43FAOtRiDRGfmCTLC1Bxtrjz
kDflwdswrQUEIGZRe9gUTyHr25TkjlOviSsKXXHYJ4H/FW1e0RZe4dzfpP+zITvi8bDA52PPa3Lo
GADhaekvnklPEcgBUuqlrL6LSNIVy/sbf1Wv3ITo+eEojB+uQtZXS1ylZU9RU6WdFV1qwFJbRO3X
w2BhwhP4mblNH9gSjmNmZw6/UODMPExubAg/XXKFaoY+n2iCnL4ZvUlkbgryvwbTGN9c2q1PN9H8
Wub6gJnBAtb901DsTb0QiCDOyqaFgHFbPp8uUGAQt2++Hq07o2rlj+wlxi0DfRo6WFsuFxVyYyc9
TfteOLQuL5eKFVR8eQqVF8q8h0QFA04qQ7duAkrZRu9NEjQB9LyK2qjLTj0KYNXhs8K+JomBx2bg
J2JOfUbb17UVEu7rrCNOiu6Buv0GrNOvTliC+WiTQleP69EQIGrjqBpFLB/UfGDIzzpDQvgNjCh+
aJUOxR+B8+iiGQ2V8YNBYsdFu52FUyDPyan7XrtMtwQgKbKWwllmTs9d+SMayX3X9zqoQFHcMs3R
Sg690y1yaMr0AVtJnby3k7rBLzgIzof5SZnyhZAwYIA36OeZuJJbo7kNVbw3Rx6iy2eCEivpYAnk
nlKhKpg9vab6CSguUiBwS6sprNMY2oDWtHhv8k4TcqM7ak+tYR8tD44ce4LPBOf6XhhB8jdsBadW
1lyWhgofMrqFSyEmqtuLOwM/kU295aAcHpdwQdjGST7mR3py0VecsQKSGqwKNVwSZvKWhRHhQpcH
fKNwLH1XkPCKPVcdKvxDaOs0cZDMaHLK5mooALRbWnQOJqcC558o37SDNcDx6SpPaILmXbgAjjEW
oAOCE+lPeV7pNAhzkDseSrJfAavrFVmln4JTjjer6bzxhe6XLY/0i2sHjkqDrq2h25wdwuV2JJLB
F74LP9gH7lv+qZEMnXJmolL4j775Z1M+M5OV1iLFV+sOKGBIBnamFxPlAax12w1Y29GlsHW4yFMz
1MQNJg6QLtdzmOnZhnXifpFuou8L+IvHW5RdJtWrxRLjIBJS5heYsNuQD85aki9OBdaFttBf/wVZ
h+Y1qwhGJ2wFW6HmIQp7fodPZ7y36tfUozBL8m+lIbHxeAqahV+Y5WuOqVqPwxUiQeibqsTNzwaY
240AlTml393LvT7S4wurdhRyIEBGjTA4ZakfqDEpM+rmI+nL75vPENxMvrUq0SMS9ogZ/V+PsjJK
+PCUEenzW2IblZbOBKi1A1HS2XA7ppGH3pzWWplWMYsp+phOtFvFJO+vDTScQ9FUE1Z+M9C1jMvD
OKOoNP0B16lXAOEpwJnBP+AMpv71ByHK2HkANNQvDmRAMde2RIbBNrQvOVzmKMDge7N/GkSw1pO5
EnVac1CugMthicHkpKW8tz8PgtV7iuFk/+tK1mbh3y1pxU6koIo/7EfpzejkOhL71z6wkl7lzlR4
iH9CX6XLFjAeEVIQajuBf7dzwQpu9dCVSirzGwrjplQ64bMAwVkQ08m/Tl3FxnnEAxQRYP6LddjW
R0QCPFQEOaZdYhj57k8s8m36s0OOrRJrB4gmZxmzqa2hiUmcnoIIkho01GcytWA/TObiSqATdGeq
nsjIV4u7aYT9Dc53BsflpMcnUrDHJKDDhEeCSLodsFch7E1m4K9ZjNLPobo6e6X89BETiHF8kXEI
kZqDpXaXDQo/pJxjwDR7dwChvM1cHki4P3trGdzUkrnIXk0833nGHov7xBP9QslY3EEq5ZXqDSsz
UtCNOqyzaK39i3+pM5jF2GNi8CwlC6szdCJImU3lrlyt2i0jwH3FmYthn3oulQW0eT8ztn1FofSR
4VyD9faImknBaHl4ItsNP9DZ8ZpVNp3jzlvxWbVkhyADoitPFDNMKDQcnIomYDrsP96Sr7vRxdbC
Z0hMOP4vQY79lKe7E+3aPkt0s1qongpjMOd6cti80YEd/z8FdyH9k0GTKqZU09LpJNsqAYxKu86c
bEzWogBeV8n3grid2O7/LOmdYEp40K66xqQAwv3G7n3ZbuMWvOeIutE5yO4QACIb3lw7y392H5Zi
dMWQ+8IQlc37ZG9Bi/KSBkeI4Hu9AxCb5FhSXUPv+JX1wnTACyS8w5NNT1WnSJjvu+QFGibsh4+2
6rQfLpcj2S6YbgyfgRME76TjrDjHawdebpheXTKq+KmIhLfMBO1m5m8keVJJoe/enyG0w/K2nsVj
Ru8G2N9b1nDw/MgtzqWCnm8tqFrlJbjQxRKWuekbA/K8sggX3GjqwUnXXswZm3RekcMcKbRw/a9m
i2mdPtjBWQd9wcgzZ+vFz6CRcrRrs1E7EjiU3ZKnAix9zQFyW/QOPFTznXcDeAbC/g0jualfToBq
y/yuFN2mZuvfBWPVO1Vb7GbSeOq85V/eWWALKKdTrMmRJzbqIJj0/KxyREB6wFUgQqVgjWjit054
l2rC736moLqEYsl5UOzoFxii66bHVMfJObXiiP4yzv/WiA9ayC8rKIC60blFdYIOCmjHhrSoqwBr
BkRR4wCwZTfygKDLzvlfI7n6d78WUq9VJYAu/PY/GenkCTW37eHGIdnwuXY2g81MG00SR/QVabP5
GcV7StMpQ3NSWzfCJjXfXR4U4cSd0qXPLIhBsOk4IMBL/1fsWqydWA7q7UTe32XU5af3ELpFQT1l
OQxEkkv+MnEXM8/yZTrYE/F8ZzNgcCPaXd0J9S4oWKu5hTTGga+Q47VnZVqQNmBeBGJG6sKsakTA
Y/LkaMb0Yx3V1oSXUR99xJcoDgr/raNhyfWyqQ5sxWXPOxr2Frne8xxiI3aK3OdRPqCbc7ZwrdYE
Tn/i8Fco2mfWGgHgedfbph9rcWaZQt8HJpD8aHXE+C7mbAX1LXAeJhteK5nlJGZHEhfMYaAHGy3s
qIsapXIFQF8L5vPixgTZuxO8i8FIAZ2pFsiexaQZXQMkeaA64G5BWRbVkPlRLJY2a++LtyUOyor5
6EUYGn5lVJYom02LPkkwoEpWGkkHzqaoS0AHTXcIwL1FPUX13rERNQk1LHgp4gL2J/UtkZM1GOMo
m0kNNWBMC3PnP7EPZgwiOWirZtBdpwjJx9cSM29k7CXkRBK8wc27HYOb6TOR/Wci20FTqtqOoM1K
gTx4ZL3ArFvhJWHxnXS7XZsYEIl+tCvrLq6CuEGuHQ7/i6616EDKqanozrseV+jwMaKjG+M/SE9I
uhsxd9El9UgV+ZlEOKJa5lWGmviF+/DT37Zz2KTEsU99KqSrJBm6kk/7BCGvZOB2k1vDD2khBhu7
NGePKDfZlLU5h8NFW41bmcTcXNw+gkFC1RWaHVpd6SeTerPRXCJNYauS7OWM9f+5FCVRWA73Cf6I
JYEyWDD2vIzeFoubAsVujpBz2iGKcYIilM1OUG+MfYqulYJMPcv7idhT0drvdoWNP5HsDSQwN+X2
9gs2KPVMcUwk1x0jTvdmrDyFOMD9mwZlq2T/DH7EmBp+zrH+1CoLoCicJueEzBFWLKwshuRktFba
XOjEYfE8QyT9f8hJyVg+JNjhjvB3mmBpp3k/JLJKVpwUahEv9L0jw0vDGsCP6bLEUEHm1kRkH+hd
/Srk8PeJsAVgHHMId/DVt7SnPCkWgVV2v0vC7uzRKZ3KTVMMqdTk7iO8cLLepUfHs1cfLttONARz
Yp5TMsQFEhc7DJYi+i/ztHcZVSb4n8I6UBtUs9cErbDJtWkVK7TDS9c27F5sMps+VLSCiPpf13Jn
lAtnWtafF/bpc/Qlif6y5KmIj73GTrOxzmU7tDIN5aJIZYFm+Ytv6xuHDgayaVfp2pY3QyVwRkdM
9aOsSbBL2yZwTrZMZZrjhNWEia4GWUui2ZiQHHXUtw7Dp1apGITNN+e4VwL4DftuEkN55xu9itfk
OtyQXUiDqk9ZTk1c9FZOirmru9y2d3A48mwU5J+xqpoScUukseGnMKzI7NK3mFQYyk0w5L4fmz4K
CUzAwYiLzM50cWUGddOWADpbCRaSi8bZZ2nEwCRvVdtKMBfAmYq9JLObzyviR4pAJP9NFoD+gaZk
YfG4E+1UwoFtUXdWiWye0FEKaZfWD7pfPWsvrzh0n8JfKk6dL1WZN+Ww6ZuJ3HEjhOEn/LIHoEq7
Vi0wyjLKtoVVvxYUsHDmct2VcF5H2kYSSpo6Mq2xPS1XlIJJVT81huckxDXsNvBzbVrWBeiaLP3z
JavqBNGyYNLdB0aqJ0ZURr+TuvRn8MyVUDsRz1sN8/nyrO73g+5JIsCvLvccn7nn1euckfcOGTtX
KPSlEr1KgNuV6MIwjRj4JKNugKZx6KjGF7HamG2jGbIqJSjKhBDaVcA8vB0LwXEaQhPP1kSI41xY
jsqtT/1zW2oPAlXjJ6qrLh5qPhOxBhWXlUApCzw+8c5kyzVt6g+cl+gJyD+mscuI6Ejeb1g1J9gL
0zp3UNzMutogMsWjGtdrqtXfBEi4rLo/qCVy0NqwUqLL2GeKWkJe0oRY/hCBj979EwYb+PptNUJ1
FuC7+Sh5MweW1mFNkzdp4jUnCzMjSc9gVPUcAHZhf37st7Qe+hLyQoL8hoOH9Iqb8CA5fnWl81zD
qKXrjQcyRxwJftn7+TOoPLkbo2PwzwlOqMz/peCk9g1bePDvvDPTtKXySJF+p9trH66BydO//0HE
jMOoq9u8xzOsQKvHQOW0LNBrp2d5cxLLOYZ1PGMOmoTyYTYCPaAy+PQUCqFCxMyWc/Txk2QddWlp
U8KkfuT+OMEry+zV1MpoxVcX2oP/yzE9L44/4T7CmfqcNx2F9VZuqq41gi/3008SyDKExoqUsixz
AIztOlDpbTyDXp0KNVEikyB+IwzFKOMyxfQZvneDtgenA0psVYUR6C8kpHbHGatUzdYzK5VhfBcU
J9gPpGcE+3XkXy3m1tXF/sDC74pzOjStq8jJhfaFDokxRC5YNDElaq9chXYJpR0GUxZ/LmFepIXo
s9aXi0fSdwfZV/Bh3TPaZyK1BPdoigFtb0+aOfd9YfR96molH7xtWtNKIL/aOo+YeyvQHlTvKgsN
S28jqq36Ras1TL5Sfo957G4cgtpTR1wzxwnLpcGQ2qRDBfMb+aVgak/hovWbBIF+VqZd0nQ144bx
0Bd+s11FS48wVc3MOIfkPsCEE62XjuUxAvTaXeOZ4d99p1d/crcfYrXZzLk/uze/OcNFyqf0r4qK
mFUUP6aDZ4d051NutDwf2/dr/UJdBz0AAH0M4qT3SqDW9zlm1onUa5pDT/Bcp51MeWSXaTBdi7E9
/ruA7ZDy5uId2RHsiJByc26Ou4mmiGt9Y0X6VdpC9ZXaJtHAhSBVqzv/4FTN3rQokjMnT2v8shzy
ilIPLGi5k1sZTjcd6FlQZUCWtNbDVa4lrug2z35N6DsPWkovEO6Xv6xgnVdSDm5UkdVbd9/zk9rU
hUpX4a84Xj3jwjx3DvbsgcYYuH4TDFs1Ym2ussS3Mty2s05YiePryUUJe/9u+WSxYkbGHPE7dRhc
Y7CUrDOCHDuAA5xzm0+/4CjBwiz2AqILUkE2qKzKbalb43nFlMM5xGbk4b2NCfno29IN/pJRPs52
VSCEzBpd4WFRL8Utf3i8E68MgW3Xg9DjGR3EhKcv90X6VCQeOG4CzkjTwSUHgsnPjFkrethgJcWC
R/XgnRhhUcbwo23NKApIpN1/165P2MCjwggT8V5CnhZx/HZucGxxaZF1kPIhp1XguUi7+YenfSzf
xnnJwAUO6lQX562CVVy/zKl3fBKJRj6mEGFOh16lD4eM0SFf96theg136wgkT0VkWMTCtY42Q1f5
ZZj/te9ihplZKOLEAVjBvkgRfqSNnRsD/DnK7l2m9d3DHGGiS71cafOdbXbVDuHv3CzhT0xlZr0a
E22LCqs/8VZCQ4Z3OpsfMvUWPCYEJcmqJuXB818VrSOTKVhKhZg0GvKrX8yqB4HwUfBY3idYgmXM
icRuKZIWlIRmVi0BExT9YWQpcbvs4JkvVKe90KWEBSzfU4Qwr+NLmPDF3y8IP3SbsEHhjv+cZk8P
O6VjTrK2uqtkV6kEGWZil0XDYzJG8M3NS9GwcfdYewuUcQlKBYHPjHj3odC7tMqbF1IiMuSA0ljz
4H0t7ZELtCI9ST/Dtqi+sRYju19ib8VtD0Z3UeQOtyJgNTI2Cc88KW+V2QAJLGOzpZVztZbTDUyb
ZcIle16dmLP1RTjeo1V2+R0QFKCkkl+A9oqL1ocUhuiIkq+ySv85ZykWxWPcjjBVIXK2OFejVuMl
Dkjvq8EQiOtrjJG0hXK9aTaEfBQIPwOAEPzTCDoC1ClshjG2yssO9IkKVSlA0pO9AvSghUK84PDL
5mKBzZeG8Iz4yV+y00wc3zxJeES3+pGK9k0+nj9JIFOu4Ca7tXA956+grBPT/MkKumb/wL2tmkHP
THBS9fDceiM+dGXUQ98ClMyhbqrJzkTSogfMrS94KwHBOSdjTs5oktC5Y7SrJPqOt5GSef6MRgT9
NsKfAPEefYaqKLQkt5oC46MKEh464GXvFeVePaHg7xsNxv3XP0YLO/aoCYPYJNZWQCpiwhsG4LXR
dpRkTuBMPRfye/d9HmvRUdnNksAV3MBOsltvo225TMQD3I03pqur4UT8NkdDcZjYCdG9ivvc75Rm
fQKDmwYv1iz1i8LXmH8NoJtr7fNujCHMcBb4hBf0jTRA/ms5FxEczZOaAnnTTK3kjQm8ru+5e5bi
lGTxIfC01+B7UX61v0b3uQgi88GCuw+E8PcUZlqHaxlJK134TXI0UrDEx2xib/gOFj+npYMomBEZ
EbVJwjIRMhwnamkG0BDc4r9lwYEugvWa0GmhNnLybiwcZA342a0Z4cZ4RbtB06kfuQM9s7MiqIvi
9bnyjSTMzovnq4pJruJHi/XM4XIc4ehEZzopAcN6uRK2+kytdMMXi3uq8qFX9mYOIiLh0hnl9cP0
xl+teLGHz6Baai3SLe60oK5qlyD+GX1hOI1uBXI101H7GcjlCoOyKQtxD9vWaXgPXmqWhNaAE0Ck
E8Yc3vyvtt2tpM62GrHrDR83f/+MDM5lWrYbnrQbQYNGYkV0YnT0djYQ6ESeeePDz0HCif3Wb3uY
xV8eWDoNOTYhw79Y0GghuhGrvngd5e+wJJVj5BzfQazopkRlwyZzX+TExyZA5vmlmKNMJKQtBoPk
Qx9IQQyD67C+GPjKfWz6EpQ9r1EEwwReLl+DO3UyRflKIEKNy7x1QGobOWwYusLynt3o1TYLlCrU
tbcn5DQUXG4mzBv5uHCnXFS7xgsj8/Sju0vrZVwcd0pEHAEz0tyDF18/S29MyvQUUVN3TqvWgOuN
m1ctpH5jEQQlLGY/OI1VGlY7qHubn9ZhescYgxZYWCRWYblgxBOavj8xMgf8jzkTw2Glhce0t38d
4N0Gu9g4EkkXGYKrhmGdcqAuFZ5tyrXaq0hZBTnh5BYlfwNBsw2Wydv13n6PzPi7VShlbN0eQdVC
CtES9CYG8CGAsyuyv6jLoMKc2TBz1ZJsm2xMlo8i4LxNHkWWFUMP9Kvc6cdbsN8M/XF+3QWC1Um9
G+pfxRjCgHb4mDmjxp2FGqaPnV6O5fy/W9Nh3oxsaPvlUfjXx3kt1UlGHkCjdlVGs6szc9afhdVB
8l0RJlB5DpmIuZT73tWkLU1iknvV+MCzJmu2ljsk6H8e7+cNs1hZpDYVFHLEKjEZUS9RykcE1KPK
9R9Ck13djOKg6hg5zya9YbfFw4+GRst+YzXfhFQaXZk9fVhpXLwrM66IJMUF1bCBTT64DSnFZXni
sA96peh84iB2B8fUzLkcMOXtyPexh3sI+c1WaUCGLn6ziec0yhkr/rIuyCLjpW2qusr6hXwn2HHx
0xDaw+Ck61At/D1nRZZYSMFWzAg6D0StFPmtvrQWn5o5+zT11SDgKkcIL4oYZJm/43oym+ND/4gD
7yfTAeYRyF5op/VPAdt5SIXRg1M+qPJ9LKdjXAOrmnCBITiQNgrnWBNx0QDe13YkxcBHDbZyD/qk
d7gzKstD5DUB8M5xsaPCRrpq2ddXqYDfzwYB3HNmykH2FO7sWqrrwSrBBseogR8fpTjQ6bErlHN8
QnCSbf3dIlyrIf1LFmDhMuSEvjpa13dfHq/cRwkzCYemL2OXbA0y3uzWmV3dEwXA5H0pTzvrEhz4
ZeGNQNJuYkMul0OhcHEK4HU7REBBgNtA8dUieN3MkKzSlIitPvuWFl4+mh0uMAkA5SrRiwYvBNyM
itZEJ1ZAqfy0HzviekqewJ8pTH6yAgyWMQbi9ePzCxNfMx9vV9LclJstlekPoAeqRM3GOj9xWdEx
XINQ0MpoBT96r3KSOWrg8jeDBv9PDkipC/bu3NDaJpvE/opdlYf6sj10dSCB2nF+pgrgQEAYRcie
ENkHhcqvXMleE7+MF0ADBm17y2P/GkSJfXtmDfe2IXIZgVqnBd1Rl0chv/Gx13Dn4GjcFwlfiSNJ
EBLaVD4dET+F/GBM0jshU7OMtR1Zs+tRanGsbbT7WyqxojTd6nvpWjrPwBt707Gna/6U05T+wJti
nR2oljuHxfI86i6Gb4GvSgvYkxBH0J5V3DpKCuqm1DSjLGG1S+9hQTLNxU9WH9NI04AB4IslcLEd
ZVMOTqLI9OmSYZ/ojNr5c0Mz902nXDo831+K4KO8GcWH4a1l4JBzsMJJGxnh9MVgCWMuTFM1V6oX
XNI/U2KPEbh6Ph80xo3L4xvhkQqguobJAycjvwm8ykuPM13QEci1ca/BBzhypy0Sh8IOr3DRgcBA
3hBxbFLSDK01js/vCXMn+Aryt6XsnCTvXgE1PlQyZBVJyHopfE62jZqtwQWokVq1zOQwDC4g6kE2
dMBb1WdKQp7hCtaOwA21MK65BN41GZv5tG1rN0phD1EEkM4dA9xAJlL9Cg/NAgTtWVzhw0Wr7eqD
DOTyz1CVJPEIILE1vV3pHqDQIBRpYGRrlh3txsCZ8uMy6lGxihJ9uXF3e5YmlgHLzqta09he/pT+
zXF9UmOcqdCEtsnnXxEPnwlg0IzPUahCaCqW2rdtlt4HdBofN6sA5H9RFHTtUYmVOkiLr48NvsVS
fnAhKE1NkJS42EuJ9JXS0iQrevuuPa8W7xAqJsq50B7qUHsNGBWVF0uQTidfB1aRvZhqoBXsvsxK
VKH+27l8rCNmMZOthG6rj/JSfdAuTKY/2Nureg19lhbrvs4sPfB7jxURfIRhNVS3xDMAjDjUSi5O
h2HO6mBa3x4A0EQmRsi/vua8nW5uoxPd48W2R7qMBq1cAatMjVMVhvwVmBWU8sE2HLbPvqX0LjIn
sRUPYddkD9vdDJbJAoKcN0Qz5RmHo9g9vFzPifiH41eMLXM8NCFwwao6XZF2ERDyOkUsQx5FpvAK
Dl1Yz2RDNf+K9PClNTuhwqFAtKEg6g23k+8NDBEXhPBPQRmD2c26lQTUgNzK0sX8CHT+4mMRhOi4
7v4ZWX0wAPbUddHqOu+AGpPFBJv1mTQk3EbVpj7p6VWbb9eEzu8IVHQAURrLbK3KopndtQfDd/mK
tuVTlD02bRIIKsjwKin65/NSddGrHu2sWfYJyyHav1Zi8QmLub6D6h0ZIPMY8tlU1OoCbU4i8kGo
+APtmbh28Us3jUtzKgfVeuinHBOx6u+/tUqRj+9ZT9cdcx6yb1mmNOvHGAI02qLyGDrL6cvS6Tyu
zi/U1DZqg5OYFD1lvowni2BCrlmCDiJC5ukAlkVLe2hWf+w2a1YArt1mHrV/BjHenzD3OjksG9y8
1AIxK4cJcDqt7U3GvRK0aljv3IPaqwQNu8qpfrJaHgj0In55VRQqFooY8aud70jpvnWvuwT4xzh9
Frtg4X6seeIYlzfsKI+KRgK/MKN6/Th95dk/igp4kqhxPjCou29TiOlPmuAbFPRgjn05SkeYNPUM
zylcuVK2Sf/6IXmSpmpRjdypR+9zSQtNSCoMc4Tf40vmkMJIzyptyDSoWScq/YTNt/LaXaaLtIJq
D1k2ds/GX7oUKK0WbkjP/Mu3Wf2TB4jjZgjGZP6EA80x8XFdgbaiXLt2PJIJJBKU5akmjM1j3C/L
puFlmLD+2HMdtDVj5/BCjt6nNzbBmLe5Z+swjHfu968yhKjM+QfPCbnUiENrK7Sp7Zy08Q8OwrgV
Y/E+my+rABqqG+IWWBUP0BJVQ4oVpV5cntARFglGFpBnKXeg+NRDXg4S0t3PXXrEtFkyTA+jMPLS
AjwiMREPUuWpKRzR0CmR1OD6CyYJ1MTONTFx4zBq1OAJKGrWllaoqo5Fz1biN6fYupIpTfxsl6Gf
/cwIQBJniVDM76XA9nUgpdc+ajosnhtlRW+q4uT+c3OpkS9aR+8rCk1edRRiiuyTg19hvo21u9Bv
NXkvKVNsAPAJUn3E5O5PQS2HTrpLa6VITRr6ofS0JuWD7FDWrUBpabBRg1ZqbMR19OdUfjDi03eM
wmV9VPPFSbqo2x3J3RP9q2p7McET+jGFC9Vb1Mc80ixGy7pW0QOYQhgVojkGR1QoBDKuyiC2T9th
hjGXgGpnn8KqabGxpuXhabWKtdVxH6EF+OMIq4CUGE+OXL5IW/i8ZycPJEu5091gkydxWeYW2OXg
5iZrkzFY/BzGfH91pOp9a1pKbQQaOEhdcQmwmxuBgFOpiIXe+qjOZLV3YpYGwpaMAgGALmxFUC3l
xv63dnJ8JyD7xfeNI8kpLI+uaMNoR0MdEkQd7QXU5+dSVjx6dVo5QjWzBNIXZCPU/4BPrqd7m/6Q
Xz7BOo163mrrM6C0uS3W9OZXIn+3UGExuE0Elaohabi9g/BA/L6YfuLpkewZiaFX9+iiBIfaLfWq
RCPW23XuNt3eWLh3vxCn+aHQuPAnOPTUnTDNh3Lu5mlSdTXUwZfMp+K7QQ64XOYGNiozfotYZEZW
Eyrhqj/rKh8ITBhSuDbWb0IYVWRC48xVQxzqNFDu+UC4xWCpi4jSVbniRRjCF+gfUU7pTzUsXT+8
4pvofhHv79mTvi9kyIxUpRT9ILA9WF6lB4hZEsK6CoWrNua/aAt23Jr3Muy+w5U9muOW6n/STok9
3YI/GCUolx1oDbE6fayhyf7naaRVYQOaX5NSQEOHbsI8jI67tu0txYfruaPeMYEC8ebjB3sFKrjA
qUa5Q5ZvKPlpGohVWUeNZX2uDjXPrM5kiNcVPcvyd2ZwKhs/pdhWI2w8QV6rB0+5nzgZ0LG40dXI
Kwp3rQYwLbiXc5gmQ+sAUS5hlHl5yz6tRaRX1ESP7D5/lH5hSQ6L8larzVUdzowb71iK2EU91Tkg
0TEQ08QEzLShs9WeLN3DPwJVmEVxMYwqHsKyclpr3gkmzu8tWWmMcG4Q4Pgscmu7VIBzHpRdJSFk
9IsGpqOQLUgJXJEmclTZj83Lvar1ul+jF+qxzQE0qBLMsp+c90d+mZirAzL9SOPQpNDe1fDy9FjV
FUUYuvAiNGbslo5hIgeYOAJKZZBuerErnB0kPx35DGM3gX7gy49ihVPepn0el1oswNJyJ3tm/P5W
d83996p59B0Jh40Ws5o++ix4QJmNS2Pz9cofDHAQNbUgqfjdJ4ty1Xd/2cUwlvR++ROeDoLpldo0
h59LwGpJnUm/ejxcu1acyK/YCymrqIM8yLgwzBMNRtmfk38LzHrTynS9DXPx0iIyQ2pAW7Wphsoe
y+V5avFQ8Phz1gNjhkO3d+DewDJuLmLvMks2afa4VYf8O2xDJFoDlfEj8gWKnB+qcNE5GRxFltXH
YkLuuqgDp0RXix9IPDOTNkEU/TVRWUmDEx3ubv0rdm/jb+TbpFl1schse5YZ4thZoIu2cicAYkV/
bstubucpuBoMzrd1U9CrjBadSw6qL7CGDozU0f51gEwcrr8e3+V6qKZiSJvmLPnh5GaYb5UunzVS
n5BL7lglGUsKJ82h+7L35spQIkgCJ/IG3gV7uIy2gnyRgTZNxdHl9U3gQoj6J4iZB8P1uV7YsipR
mrMuqj120SUrXyMQ3O51m6wasNYYRn9QrWlMR9+9dWAZxxV8hDEAB1cPZpIfOSuaFvJfWLNY97fm
AYqzWUwOEwXP3r6Edk5VljRQ/mv16q6T/lDt6yG8a0XRWcvw9tIdWHdgbeNmXGYX21HfFob/w+b3
QN6wSsuQjjCi6bpTut2B+Aq3Hp6LG7hTw9RBGdT765RyL+K/2yw60kXVsDU8Kkoo+hR2Q1v4vjwg
aGepKB2XRma7LgsV57hGjGq5SUaRbLBr/CfEkwAxfnE1PFuMsmO9SmioSJxPURNvQq585yu1h8op
P+PI1jd0MsGGa1e3e2T8dZCV7C2bOyxCd2J6qk2ZVxYot6W5SF9veH+M+VP2BQKeGxPZX6IH30Bs
7AA9HQrQig8D4UhjMmoLhqIUiTfO5NMPZ/FzA5aiYMaEUG3GcQfnFs0skrlSAxzQKXqDnvRTVI5A
qX76ByICuF0y9sjTRgu2cLwn3Bah5smPk+RogPusbJMcaoLEAYOT9e5T4U/0V1dvshPUjgSBlztN
4OXX2G2WtiFhIUynPOdITJNabgdLlLi5bylQfzwB94rdZ0jyrjbMVhvfpD1onVy8/6LdZVOoejx+
YY95S5da+ufd1+WH6y1ljqcrlG2nm8HUhHDSUZ+r/flAuGw0MqVrvT2c09WQWBRis+/WK0iut/4Q
EdHQ/ajrUdg02exyAdK/81soh7cartpEaQMeER0UVWQmZcYV9W4150LhDGJh4f1BAl+GcxIMm0lP
2pl3IIZYJ13YB5+HGXVknREzBs3Ru8lN6sNe1mXTWD9lt5RfqdXBXzlfpfo2VMFPH8OeCxJ7iY9+
H77btwaiXEkF+4KOcGoetarnFhuoyH2B1oqpe6/zslc2lt9/WSV0RauRfBZsr133FWQXgqjNwPGS
Exmq0nBb5brb6zBlzIGOBGnXgupdREF5oP0YcMsuN2e7X4sF0AwxBcQL3zGBoybbV4v4GthJU2Qc
jBYmzz/WXeORzEWHlS4fjDihsmRUAnhPDyumUh9pyoeqBLHHfSMFDnOY8FcyL9lht81qwGxSg89c
CYt00/tH6Zy8C4gz2N8qus7Tvj8SxE3T+mrz0XAuP4XW++lH7AN4tN87ocJeh0ETwc+THbOzDHNw
vjj05vEpmRJTHGjm8uevHN/zQwUTfZyvJZNaORLG4q+Gi3OpJpzNKg1uH2THQ244qAkEHxj7q3LT
u0xGVKCuGf2KovhYCQFuy5Gr0FtuxXICG455D1W732VvZBj5UldPfGdTyGn753VzPConixoqhWsJ
m1PDg+W78A34B3duHfg2HQ8+Ojpuy5Mk4xd1aSjrkDhgXjFKwNk3ALVmZfWWvhU6Flsj89mvztsY
UfGcOYJj+GQLbxMe6SM4hJIbTlt+ZJHeNpwJ9/QQOfUWDNzuxdh6I4a+ATCjuMPhTbQp4KE+EiDs
EDqunXmg8KhCyrHfGxEARe0ErMGh60jb8aokahd+1QaIZecw2JAyYcni5D+hXLugDPkxS3AL9qyZ
F+/9npy7KW3VnrRQf2xSpkmFOuWWZcXVXrWY7N3NwnIpN/3Ud0EyMBwPbTpwshGtvjY6xmcqn8kn
pMPFz3/KRNiV9+7wYhefeif7CxDrWBzvf587Y5VjPhtaW+r7jc83NTtC5aoCaWOJ66tlOhry8uIr
xgdYU6w28pNLXCaJDvQKvL8A0Ri2G9E4ykHneEdfx5LYYdkJ9wzc3lhFovuymt1CVtFvmTgKQoDI
ja9hQWdOaSWrKxA03Tb8OlKeD9nDXHhqAbuReShbkr0Ca+oOQAOpHtWH0bh4e0M2S8eJ+WxcnwAB
6EUGJzNcWX8xe92sRJqtG8oCcJ6npode/vfzTptjUoq5SBB6zhZt/Jkwm1FgDzzRFeP/JAbTSUEo
Xld+Y2J3XJk4HT9gttVnVtucFLwijZ5oxGb1JFCg7SqIfJlRkUOijDUqkJLwACjh+gROG29ZGqE1
Y6owUzc9VaKwEjP82pxKrVIzD0i6rUT7ym9lrbodoY++FBWHlCvRstIYigWT7R+SspKszDsSeEWy
+zUGGb4LoL1+NpCWRC9A6RGw9YmtIyMN6abU30bCUZB4+JqSEoGPHU2Re7wiEOMyFdp7iHxfuIEc
yA1qbWw/d2tAKBIdH8QZXS/gFUinyXv2FLFCKcBAJzJgcLZiNZ+ilvPc42jyKWYcr03pUWHyHZ5i
d+UH/DxPmDA4cITbrdFtJ+4ANeXFODeyLOt/fJxV3W2HJ5uvD7zsTTuMgzcrQbPXvNcj7Gwb+tbo
oZicyp6bDCIvUopVNyK6xLbcmjk8bYL6W8dlWx66k3EA5Ez8xBfBTqKuRdAhDhDxlRSNbKaKGACg
DgsNYswfoctpwc361od+ABhil1YNJmadeczfNoVBeV7lMmZ+0YrvZUo+mxFAzA0gHKUD/QlaM1aO
tgSSB8znz9JwvnXmWUgkel2Yw7+SZgSOMG1IuoB3jH6H8sGvDye/a7R5EkYKrcLhMP6lC58vBLqB
iuj93RIIg3mxH3epeX/GTfoOHrp0M+XJEsoNjBuO3VG8X5dA0m2ovM9zWYmXqEAJLNGDjN80tG9R
l+A2TCPixSjfJcS2Uo7s32txANkZq4tcdo1jGrLlHSUSVlBISXblwWr/kugVtEKJQv2AlyVwslD3
4R9ORT3JGdveDZMF8fDXlECnymNj2bj7y6RxOu30Y0+FSx2idj8zc5FHna8bmYreits03htIjdFQ
AkYRFoJ7C9NjKLqjSsW0hcIOV3ExknhTXvI7vdX/CrEkbL6WwD+euTJ6BwSs9I2KHq9Nn/DJrBpd
f7NQEXfpgJ4C+uA7rRgbDhZ09CyaWxuHMuptgdOixoODZ+ZRsfcskAB9H5+uNR7aCdO8XcDNzj3J
kHbr1MOY/me5IZhVCYu4/IjcwQRz3MLT4lnxIIwj+7+faimCaLEYSsinJ/hHWltsYuot7Ulka6BJ
HdhmeANgPZrYuq7Rf8Rn/U+bfydBWR/KBwLTl90g9sk0YtmtPAGDAQenRUqfRYBcKpTb7r9938Pb
K400YUFrOi6DYoSaSEdaKHogl3nqspP+Q3dpV8wFBc8VYRNEozQ3aIXe/puU7F0t9TMf3bx7txsA
2rhptjCu6TadBjRavAAK19DzztOrbu91Ce0L9WE0pgiF73DHzY76SPCCI1B/J3IoZ9iCstRlxBgY
iJz//+Hxhngj23If0kWi+dXVolGRTFIRnLkuSjH4SVXEAnLRXDcrfW3+J4pYVbr+Ahzh/0V/JSYc
QTU0rSjME8UKlQu7pRjmsqrDX969ZNceRLxtJ1ZA51/R5NQ8LUmKvPp4lMVNzmTkxgwfPTQFMFyr
YdJOc4j1vXEB7ostwPG8G+LL8sc9lbjV1Eqf4YuzD11mQSBzJn+1GgDOuIFYkpxARq58TjMzDjHA
btms3i8XTcWcaS874hOk1atSyPv0UWPCp4ixU00+lr8kaUJql1+EJGa28YR06M8HUntfCKdC8CEf
0grK+3BhvOJaDukEcEgS1bXpG37FKpfbZbUO4Kr1ISMu0dd4gJpMU9YwYSgt8IzCnjkB91C94kGY
pnE9aIe38gyINbOmXqfHzQPCF9tCYNcMcOAA7t5c3NJeeTUMx88KFo9qhKCEV51EwU9lPApvc0fV
WAJDidPuWSKU/TUofihhB9S7JoPCBrX9Zu2uCuKxnNixtGdBUufg4eh0p9S6cRHBdPDo4rNd2iUT
XgvNainwSEqnGsm3YtitdlA704MtM1/DyBzpu1F8N4n+7bbqK5KGHr7Ol9J1meFTbCao6Ibv6dw6
/SRve4VGyyP7WEGEJQk1tmUQh23DKa6qCZ1BA9YFj514QbINUna5LD9TLhxCN7HmFfhSG4kKshxv
CLT2YYEMFTr4NNuLLDgoug+izupiBYeN0TfHw4WZJwdXBI6cOpK8h0EhMupgm4hl8VehonE/hdRd
hADrYOkcEcybJrMeqIKI1bHgbZ5YbCUpOvp9rH2JHBB4Qs/rhfahQLC6JuUfEgBB82nSiawJ8Vm4
xWiIJSkXXALAQDiSzXshjSfKDXfBxXJBM3FE5LrfXZgcoJEo7VcIgB/K6rGf5NCGZycmB3Fli/Ba
avR2XmBjg3TPsk6P6hhHCnL4//G2Z0bqLG45mbDmd4Ov3PP4Y9+ev43mdzzgPs6jdf1B3zoHtk6d
MyLJEA3GIblghF2NHX1deen+En/vU6RTS0QfJ2m05uMajIVEVjAj3tUKZhdPF3BofQModEm1ahdq
NxIaO1z3vwDDsIqKuS2LXW8qONpvdp2GFwleYrSh7kpgFk+F2BA4hbMqeIpjFlJvUgwePB+NuGcC
dwnpIgPIBW8KKybly7uUe1f3+b8KKtMGw632SeUJ5RrQGpe+JHTGkmhz5RSKP13NhciQ/M4OHfvE
vo2C4Mpocc6F9uSsr+8mtSg5K7G36MI9zZhHpti2duCUHxplQxMRW0gZUQn46xm9QY008bE5Z9Eg
NPz31NVlupTZRr654hrpNxYLT66v5X6X2Sei9SlmbRY43W8cUQ8A6jXHsMjIcm5WJgzOrCB+0knx
PV80IZCqY0XAZvTj0axtmP4nBqD8NgXn93ML7y0sEnGYonC6on1jMhYhvmkY92yF2gx9/D6h6Zm3
NqGhdMwvhvW4OOrQL520fyLIlTdVOh5cEShAK2GNh9wZf46l9nK8TeieellEPjWJAhX4bVS45lVN
u9Awu4svkZCWSnmKSkHafDDDzHYkIb/yoEP+/QOkPx8XcE3Jn8j7eLwBq8OomHRMLBHPS5G+MpDh
wdu7IiqmLYmJdlc52doeySN3tExKEqWQXxtiZwWglZ4W9nJbx8LANzTZc++AMgkLeLhOIVLFeW4J
5Z/iHy8mql1QPTcWqjPiT4BH0PBQbuVHOhJJCkyDc75dlgDhLfd0KAdFlxka7ZcdPMQDUg0ofyVO
ptcokrYQbFOnMsziAgFAXBLKYq8+B3FnAvU4IXLud/0JuGyR71+RKqQug3RG/vC30vaaMsNT75Y2
Z0g14EP9zmx9aptYA/BcBnbuGtrigj4PjqAEwlxere3fiA6fGiMMdfOs6vI8MuOF8xqMsTXGqpnA
87M8qK3FTwVz1H99MuQiMvJRxCaWp6AoYcl2kr465s/pkKn0JkyIQK8v0Hgiv7GSo4EfZCKtjlkU
ga7WbA4lCt7JT87W1b2kMarkndo1krIHC6jdY2JnnEXVcL5qXTGQD1KpyBSbSAC5MW/9Pz2jrzG8
OQpSOT0mAxGL2JOuv8B6x7owHk3gL1sWjO4n0zPUOtqWdT2y77KqGA5/0s0/86YI4w7mo4TIjMbR
4DaKDu0ot2+47MicEpeycqUavdqzM24Vtm/OTIsrwbGBZOQoCOKgk+U0uGlG3/cfXlelD/So+/D4
J/ypCYpXyU+NlRPVdU7yhsLklankEw7USy5761wsFYtejDTU6bk4ZRmSMH7QaEAKPxpYqn1MNV9O
KDEpwatoN+QXgHXTucMH3dTV2ovUuvZIGKmlQuCpbEg0RuqTIN6tebc6uiYT2oW9QLMhe9DhukQo
9D0AnXWqgvrEhMO/VE5wRaElQ0Yo/cmf2pLkjwPqgzKyNgq/0BUrFHgjQlnG9ko45SaQ9r/YLEC5
QKkz4iEvAYHfyNca719Y0D3ozgeCI9MoalhEJhhKqdTiVyLFcJdN7Xl32gPe7WEGtvaZOTGKdcTS
Yz+iMHZTaY2Nl1kWBOx8Y9yPk6KYK88nyEkxKwYtY8dM4+/XP8e38TMB+wEwxc65g8TfhlTsmyrm
yWXk02vFknEG7ymP3Qd7GiYBNk1Cogk/J2uP049SU88Yg5I7uSWMgk6UIMY8ooGhsTmmNjiHF2cP
clTg0TPtTKgTGLbA68WRvAyXcgK46XanYtEN6lTGQx6wkAFhYOkm+cZ/MkhuTfIL6JmTIEqA0LQj
nHq9U3RH6tu7jGdmL4Ogvtsobg3Wz/r8+hPJvxPnxSfgq0NOz55tp7sqTQF+knPN0g6tJQ2h22gm
egAnhp1aqh4NUwZbDSnt2ZuTlmeERdVy2GoaWlcvgaagyOa2w68qQSNr0XT0eS+2tAX78n3puiy1
LphUf99UGhoD+/JVcgkSy8c5aYK9DyqgIvlADTR5VRZ7T0oLE2OKv4MrsBykvlb7P7P472P2R77m
BiK8KKx1TuixAXQGMLC2+I1Ih8uAHcNTIN+cZEfJx6MtIi2pkfHgjC4YAcMorpCDTxrTFjwDFkOJ
ulXQOyAOveYpPJ8MbJ0aX83M+/SZSxxdLtdIHxdXh+4I92W+7RWILDfbVMPidGg7Pa/93Ohe8ff3
2MW6J3Yz/i2SvF8QU3gNw+vShFksMhM7GqhxiXGeQgqG8YSoVr9RThHq85uPll4un6UiTJKMl5lL
3nT4+yiQHO+OtbmiudHoCUYccu5gtPsNZUnKW+SybfIN2MRGa4bWv7nJpk19qpbIQ+AA2JWKv4KP
WJSfplAhCRbcTXKi0XVZUsQiLDdYx53GP+cj2Ae4UANa0mAZIEYLJCTGPqg6yrDGglXJFGGriKu+
hPGnX8Z5EES2J2XoZLH7V4QKqHRl+iK6IDdtGo/cPW1ZVM4n7bZYIrAL2sFSG6ZenRMYI1Wnr70e
n76CLVsqf8U7G4W2p1GGE8rfks0AdvVmWVp+iTKD+Uwefgmbj7uAgQMR8b3zVPZP7lqtwMYeMd44
+1BAiWwKktNB+1QARNLhryXqI802s4D+KR9a2bfEqRU4IM/SHrM9JaxTAqLp3GiwfVxgxwKjLFfb
mLv5xpDBGNmpY73rJBvEfqqB6QRJTVID6usBgJxr7wyqmRDRhnuRGZNM7NFhXHXmt8c/t66r4+/Z
RqCGF84NZ/bYFOdaULkQ1QyvDww+idSofy6DTOjxcVmbqlcDcZHW5CGwadb19vE31KI8WCGH6yGF
e38DA5HrIs0/2G10ESTNmdTOj7NUc3ohLX1A13I3F+hnKQ2V8210NEP3Y+xUIRYZSeRqHRQsoDcn
H6qlX0YX5aFB9bZD2iObkhhJaU0898JsbUxZEx+rQsOo/F868k3gTf+3pc8djJnoQsPcZw/txtEf
oupsxM2VIN68ryjCXQD50h122Ifc1GB/MT7O0V0ZmLRjeDAi8Zivq/9vHMAdIIzLXv+dF7OjJG4i
miZpZnMTbWeDiRRweBWWSsZuV8z0JJy9PAtLiA4JR38s50MXtCbbbN59JAalxlC+p1u0cQ+i5qnn
OqbDI9axZKlJMFX67O5Y3o8gJEWADVAzLht4pTOzsm2MQlYRqPg1IqJ90PIq18o4YmKsygsRMImP
ZXophJRXbRM0A0dbj+QChJbQGKxnkLYGNE8sQEGypzzQiTG/TosCLql1sPccrAjBtBKMKyVzqi4S
wf2F8nQ4K59DLw97Fe7HHyB8kUBps8MPmhdKeuJDiFLXKEeP9TBDDLI/S2dowHiNpPFcz4kwh+yQ
MbXk3xD+4q1hU3pGua9rxGdq2Gp1KokdOjFnRi42uYSr7afW7bJocIbj77+vaGZ33TiXaiVmqDOQ
ftiddPI7XMnaOdY9HMZgOqI3NfnI1BYqWpU35DSyz7AIrYt0uhPXXn4PGQaK8yC/V2KiAN1vPFij
m2Oii3WRFQcmYDI5Nv/KeuI2E4iHsxdhTWA5CVBfBQ5Pv6xoGxzFKSd2pl13mWdnQZBMA7MVZNQi
iYKSCkD93eQsJ3VgkYEywdKXjlisXqo8i+rH6M4bwCjCXIDscXh0YYjIeQsZ7r2jODF1MYSpHIGj
8wwYFHUaktBVfUGAwzR784YQ8ieDxb8v64oeBFU6jOvfXOTMCKFY8OpEILLEsqLi7pkJ5javM1Mg
bWkErPnUAOOnmYbtDhtJq0mlCXAqZ+sZErsBrJvo499aKFDNgcbbPjZiHb8q4mVIVWYEusjDVBgl
kvjQS8aI9N5PAGH/r/GGJAqtN7okIcw8a7FYNmJCWi4N5VpMNHcPHjMDoc04Spoi+PzhEfX9Phur
BimApQg+jL5LM9M08d/fvA8deuxZwNQj3nir8ov6e6hLin3SJS0bvexW2otupMPnH98pW6gl0rKG
Uovb9wA8Cjausi6sCPjmSgeEYFp8np9TWNIL75Hw8iNTKL9qJ5QVFnQ8x6uRo8OoZlyM2MSoBuQ5
HQv1rbjMf/1ZYYytHegcqsodhY4NN5h6ZrjntdEEZIhqByz8T0cta2mQqX3LOzrJHCmPscKZ/yuD
P1d8VXT/KrBNlDdbdL1XOSYE/qYl3tH/w6aTnUh1A79kbzEL7qDG75Qm/Ma/EqR33nUTiUCRM1/r
92f6P8l+h2tiGuZF0ZWFYSVxdup3s7iwoz5TYAw1jzhP71usXIu8ensAA4ScNGBzDkrORQ8WblQd
zaw3AgMjaDEysQ1OVX4TwD5vBbQBnRwZ/GDJYGkkaxfHWvBqOlrE2+czg0vV1UvkJu+Pu8Yh2UpL
iWNChLhejGnJtMr0viY905vTXfEApSXEBggtCrH3mlLKoU7P1xiQzRmvnifuAviuNv2wPIojE1rY
wVsNprYbbe54xOi0pM3/hk2LTJiEPz/DojdT8tFxGutpVTrzvscEBtnliGfqpPyhm7NGOWCnehzJ
/d9vlYj4xP1IH7k+myG+oY5Bv2rLYFxOuBiA7GYp7p2Rnds+jp8PPsrIgZAl7raGDED1trx3Dsg4
v7LT17YeGxFmnKCzIcUCcglBDcDyC3C6DZjepOYO6AspPgST4oRLZGXCQO+1SSgcV6aI0tHUOY+J
5gPfXj6ww4DUfNJU/EdbE7/WHQbKxIw/kevQmy1VSIx++YHONzUyXLH7vlnZmdEiaFVOA4JgjNzU
vKXV4cvwsrlOPT/PXAWnjpoARy8tazzOEeGZQUyCbhG5MpAReafFHEAUhN+Rq1qCjtgq88I/hYmN
3/lLkO/LDgsnJWS9wo4xg9ZksrC68IcvIfiAEihEdpGb9Qd69mbSnRItlO5F7DigxFjEHDqSt9Wi
4xqnzMBZAP2rm0q2F0QIDFDqF+k4hg0pwAmanSahzlVhc3nqH+nEIgbJLA/2UNwYiKtQCdnZRQyD
xEzVTHt05Xsu2TOgs5t1qJEY02/8tvIUFUWc01M/3VqK5SxaBjWch4q5xjZ76ZelCx1YULGWNQcW
NNcNTZt3kMBQr54h5zeJCRWyOLDJxy67dpepigTHGqDIIqX2lwHHlsmDR8V/szT85qnEbgnp7QWh
fmgm7XCPc2GKfOS3U2kCFpQrEWiAxzKyDEXOF3G83Fs57gmG+UErAWanBg1pnJzC3IAFpqLUATZK
A7QjdlMAXRQzlf6wJ+rIWy1EcgeqwdI7mn/YiWzQeyv0eVFCOhlSwX2RjzvBQPwr9bGDWoqbW2g5
BRSKm8rC3oN+r7IWbxzIE9R7kt9Z9kltnhKlMkq8nxvEcjLT0zT/vrzUZgK2faSuI7eB8LRkl6tZ
T4CZtKVvAcoCgCdN7dXEon60pPAs9sxLhY8YJxeZ3uCleBFsFUgfHopbJQpA6s7u8Q4X8/DRfpEn
NGB7uvrG9o2SHsEBSxMt10gaISWhUlfqslJyiukXX2aYU7fBD8gVfYiLTeyrdHydC9hlVfMnGQyx
8xo3llAPOFEjqQ7+D66E6kdjpTBNdQf7FwJsK7DmZwMpfeL1FJI+D014FSNLEkX2JaJoSwyL1LJl
7FPv/rxc5VKCDqiSczfXzuSlbM9sIvqvo30UXX0x8AP46QpLEgXWZVQiwakZdobi6QR3nSOw1yli
eWVTO28NkciU1TLy/4jwvRFDMIwAw1th6RdQRftJd+Pxj1a+hnCmx/hZHtWZU38P7ed7BnhbIjiY
g2YmQItpUxHLySmgVoWblp6f/C+pyeOpvP9ByDtw2aX65p9oTwiSpyfIBuU2OdQRYKVflASYOhZA
fvfoQZw5YDF9Ri53uGvvTYPfk0uuFIZVLuRtA2q+raNhGmzz9Mo2aj+P+X6PXxpbDZIohmP5cdee
N8+f17ECE8jovF+8opGtxfbZa5YRJjkzmxBRPA1SRv0grJTy/q62Rma1fbHkNwu5uAPF19YmaLbk
E9DIJuDPTnrxNsmNDtsjUw1n73DJKRQvPSJ+q5czDcadd7zTMBgwopBwULMll52MpL7Mn//6ag+5
oIhU4RX0W5R9wDFh2/vvySQOQX1JCTTWE+QATI5UrZ4GHBtohdHIrZQ2uN3vU+vOOJwV9B8mPDIR
h9Do3iPQVgwjCV7XkMDQG7tAOFspT1iwCpWCNXFimm9f/v5SMH1oXMcIqBVafKiu39Y3hmSQ9YeG
Pjqb84LteS9hD/lnhUOA0WF8ddGGFPUKL/CjYOPCKQg9u42A2aiCGeZQKADHNva2bZ1NUDQBo77o
gZVJxxj7vy3ouNoyVgsIoE1BboYyK5MpWG+4unRQ4ijdnnKoNwmVh0GB7fVmxKEAvADdtntBJfAx
vTZ/i9/+w6WG+6oNuf/Ujbl3BdvhmGwwrbKhPPy076jAKkHfZF9at/9e7xc8QEvowHGb8iX96Ed2
KQQYzA4gZGEQCHX/ezKfjr3aS0RqglV3+QXqeYskUQa1a0KdIjuSUpC2IL669tXQ0m3LFgj/WIq9
YZCYI7C2xf8/TY+Vhpn27ZRR/T+KxvoIarph+KyhvxJ5Ih3ICGwtHVYhThtWVKp9E2lv4cCHEpbD
sESWeQnWvzHSWTjp7XoqKyozbExmW/gOMEp4ZOpVobwt+46GXch7pkn6KLXtrSDFP1vkODepN4bC
3iyLoi4zGozsm+8I/qWuM7P+lk3tZLSN7KaaatgLoPbmqIjXxWOvTtEqZ67NxDECG7P8Pu7BSdjI
XfbZGFtniVCSfOMsuQVsiR3REXgRUYdBzRoOFwWY0745E5vCoVObx5Ts8xtlbVmniq4x4GKx1ICw
RgIhqONzNMrIvAkq4IxLyF/Mt8ScHEdWhTRunRqmjBmzHBajSC8h004RPTG1PHINk8uIZp7Y2T13
Y0AQ660rITe4Dp8xetkEs5ebJkbIlU7rmIKrejxCyUkeo72Y5SOXklmhNIBSt8RneM2NnvN1f0Ys
GAZqeUJyICPqr5bOkXgLdlZymiGIsELPHDshlP4RuZ0OF4lVwaPVPRa2A1CnbW8z92+PJAnGNzW7
T0Zni+UuAY5Vq0acMQELwuSP+BaTzP2WrrDYCPXrJLdWUnq83wchQ8kjZ+kMEcbI4ogS2Df+S0Ws
VpjSkqq/xHtr79WPsDgVmdfl3poUdUjKAshyDzy9RLMsG1/KId8fNZRn+2FPM/Pa2tw5W+CBe55a
NJZbimxs2rObINgQcRLa2fCut5JUX+QG/z1fvP8ZyXAefPbhmQDcEkehhw1vF43CFoSp+rdYDijv
PefNm9jb5BHf2q/GHe3W+LArbTpSxH6auZbirBuaPmSR/cb7DlTX4pKeDoEkhcDmmq6s05WdiXot
5xwxUBjvOJ3jBJhwOwVcULw9TfGriOZSZ/oa71Bp2lj7vrNrvtZBHeZ9IY6xijixevudrDhz4Lmy
aMreMdzmUFZAJ4CMkQ19UeKk8mG6zTSzHkkVZoCd2wnU49N9A41ZRohwXnbcgzmGQxjxrL7xG/Qa
ovaddahxcQK4SbijaF5c+HoOI5DhGpz47/nOuB60QwoahZV12u5JGPw8m62XQVm+xOwBsj/Hd8/l
ml8+524H7jidZT7mLlFu1NS/L9KAkY2LVidWnYPWFxnyaaeFrZWqzLDME0ZTB6mJGP+e9dAPX0wh
DbhHNmqYLOewBG+8i5BfEM5aDCY1MSTB4pGkrXF28XkJhY0+M519sYif0zTF5D3fSLMmEfWLFPQX
WT6Cw3YSteOL5+efCz7uvQDlO9XAz3pZPUdp8zHiYL91yavme+wRv/+bgjaSeSJO27oeIPLIoxWg
9jgJhhDAEu9lkPU+/brww6nytuTDfdagC5aYDjQn4fpMQeAAq3vaU0FQHxxhU0o16xmyqO710a3I
x3toTMxzgE3DFAfx0fp2VPQpU96Tu/s+5ngcbtqXmq8qgIO2lGLXb3O7RhvR4eG6UCy3WEvF4KVL
u4+iA4Y3uNlfzlPD67f9bcH+I7Vox4a0UNY2Qf35ZeC08oLhqHVRNLj0YobKa/4XSgke5H8nhC7D
24kwWNdfCeLJvDQNqeC0dNynP4n424J3xStYjynZgvmaTVnJGm89gdZQH/RnXG+x3QLo2prbga2U
/JYAKTOAbzOOAN+P9EV6FYNiD/ikisA5ZrZEbvzOmWTN3XASIMKvSDSnBpnvgO6Jtp2NTBItKq+5
jEcf4qeG9vGJ5gqseJNUNAgIxTBuQ01Nqr8BSjpRfE2/VyQli1UHOt8kwgRiJG0PIQAtMqMxIK8T
GjJTwr7iog5izVAsy8sRoD6NCtPyBBegd1p5mhOqawbk172PYC8GNLPKXrwhN8OeC17bkBiIwcy5
5N/j+Xb2LC7IbXEofIUCq7XpRCA4eDmIZAuVJ8VBc27j9IN4eWjxT7zjicXq06OFyCBg2z8WbLV6
cCWB8ypj8Va9l6vtsm7Ski5r5nvVapFiScVXzqVFLdbJtoEu/CkpWpcn25+9nfGIwbFTdOVWpyNa
sCZwUcXBPE9Ho9fgZQ1Rn5hmCl+Q5ihBRrC+9E+uqgV6U9apH7cUWatTH/41JC6e0Vw2a7DQeKs2
g3erAy3XFCoctQMQx/Vp11GDTI186zX4gM7jzFITYdW8RQS7zt/9TQdGwKTrwRamp9x3GMASE9z3
8HxtyV1u1Uihl4YTmRGoi4dJVXtbviAM8VHxgqrOSg+lmcRbFxB+o3O8mDje4lrxUGIen6wMad9O
2MDLTjytWXGMwxT1otwM9o0m3pqUSBi7S6Z0vEEmwyhE29krE+eGgnoOas3dBr/aLasef10FHhLB
to9Gy2JL9Yv0ZqXxGVRlsPJH8ohhV9liyJ79XrWENP9O8oSs9nZuPOUP8PBafd6BoOzONcHyFvOR
tEMerlv3s3XWO86TDAE1QTzt3GN9qd/UWDbV2xfKU3q1moosgHDCQn/E4TbFw4dSxHQy6pSZWlOx
yG8+/VgaUfzbyBvVNDyhVj69uYBGoE4Z1YA/lYkWUXGlneU4ZETSdEV2n3k8vNIQ82Pgkhkpr2mA
MZv1n/sysWZfpqfygvZ4T9WSdO1MAAOPuPIUut5LBherSPkdE++E5xo2WviC1S88Iozb2PPJFv5l
Ln7T0TCHttpF9Mz4bKjfniJfDFLIRL809I1TVuF044ZhJ/m5uUKjzw1MFy2ikUA3P4xGb5X2zBXU
dXVZWvS/2AizJEiUA+Qxx+EmFMRoDK+Omi4YUxl8lnrKvxO1eeOwQcCnkuRQ8JxwuBg2VRTwXYuh
rwh+9Mwqjk0MfH5RjxX3r1eOG9peBVtEOVpaePq1y8lwrPExTTObzl0gbq+36b+o63pgW6qCPhDX
qcFx4FLCMvMC9pcJa49BVGj2iVUbi5VmKuhPrUTaMuuX4aU0ya68bMCQVavp4nA6bW4TxWo/SwIT
thiakACnSWqDH0rtWARvBn95myxj9qOi2Z5iW4TD9z7nk7wgl1GNtEBsQTqL4y1cxHjO6cd0LcEU
5es4baFxMQ+wFwKgriUTAYKdPXSy+w4D45k0Qid5myqvqGgdKMRAkvuXg2cFDf0hQS/WhS4pdEhC
0kfR+N7ysdVjY7FHfzdm20FIGXBBFV44oCboQGdXmav+w+aaKi86VpT1Of+WvU3BZQCWe5KEClHT
X9tYH6wZ6p4H/P/4dt/NdN8oyYdVvRI/C/aT3P2Qie13SydwWiNtmt3Qq0tQnIbbVPV93DofmK7I
ghIF+3kRsQ8EO03Pnrgt55TNYVaKknyHGCz2cGT09FTMe/FTXxcNjyVHkULZ7117V+L9MPbjT5fV
r3zB54be+cnQF0QrEUD6IJPySWVJoq0x6BT7lIV/sFeiHc6MzSKcON/E4NG+LC9yLZ01GUYXr0FA
F8t0iOx5H7ERx9/fznnGNR/PJYUVUOQYyHFY6E7uS8r8Ki/Zv2ZDcQZZg6A9qtHtcOgJVOZ8r5H1
MCwS4/YAmaiXCOtIbfREMS6mGXLSuCCfp1F//wMH62kinfhViBqLJ8vNHQYecfUN2N6mkncPUxh5
METnuINZXnvgqGNbENdovnrJ0H1q5+MHgeAfVDI1fRdslgSbD56HbBFHxXU9zBAO7fXBulJ8G+ec
dj4es2pFka6d4+scPU3wJfMuxrPsXgM8eZ+43a274hvOSOaNWPOcybCFBNIyq98ZNwTDS1vjYpIT
A92wxFWWg9qqvHkz7i9Szu2X+4d6zs2qrKmFSm5vNjYbeIjj+Bix2ghZlJtKFa5clGMh1WLNDnWx
zDFFQviUdlXQOEruWdqfn1rWVX0aJ0vB+OEwPbN/HPklksrF2eYnOssos3JRCIS3p/YK1HegZ+vH
8JW5YSwjG7C08WHEP/f2/hdxjvjd7yaMd5l1kw+zfktiL10OqfitGvH5RTex/hEfS1rUTVzl0eqV
b9EjxXIiyR+OjsRetQfVoATtaRBek+2j0ImaChPvpinyKxFV5ge+VOvGVXNnlNwRX9BNjtUcHc3r
haASp6a8yjM+cPi9yV5pqQyxWfhwmrSnDzDIyXVMGykNQxBR0AAVX4R+JACFFbCdvGExNN+3UyLx
xhmwglx5F7MDaRBDRj/M0I7aOSZQS8VMwv5rSA/kfRsXk9E7pZ5QHT4LjHyemHOVCQs6/43D8mek
uwCRbaFZxlf+VED/nEBXoI4LUP0wJOn2IvmieQgcU6Gq3dXYX1/9AkRZObls1o13CGqjahcgePYX
ZTFL0TyEbuFw6BzFG7e9pF+mYMJt3AlAkOlt63Odt++LhuzE/knSIbWDuYGvkTtv58NdhG1NSaim
AkeZoyW/ewMl6ROLq+v2nKdsZi+5BQKJItvUAO/0Lq0Wxmo9Q8FybaSo9UZF4h10aNaOO3vn4K2F
5HLaOSdmFQQoRiuOlnbgg3GkWKmPTX/veQ+Lwp0PhX0akX2106LmwMjcb0v6XKtUhXLs2p2jcnY6
jwX139qbZwRmMlwv7Qac+Kdl5lktAuOz+tV6Z0gccKthm6gx0v83+VNj7PbzLUPgXq8iucp2hemQ
+Vif8HTPgECZYiHjodMB88Ddum12Fi8N1vh4YLE5NqOZU+Kt3budAwrCD8xKT6LNTe+sxBwE6fNW
QAp4M6rz6I7ZiRMePUnElI+CqhlGoydrDJ5MIbz8khfb57drOrhcMH76XYr38PwtIxeRkrYU3C2K
Ndgx2biFRHbrSBc23yc9PwKvSq55dFzToF3bl36pJnQkgKoTMpKn/V4aq0rkB9M3ery6qMGldcUO
7ExpI3G2JF5TTIOeEBDSFRQ/spNcO7Uv12C3WiFQMwrUo49oOVQusv33t4CTIZCH2WSY75LKjv1I
kLmGgrrL/0WP67IiIwbHwNwV1iryXeRLq0d/iS5tMf0lVqMUgfNqXeZ7ZT0WFGQSGVghLMo7IYtE
FGxQfzMLt2L/ZVbpyUxWSTmxrfUsgcvaUKeoFdATpKOhYyMperrpxxe+oiC0fgbPZgo9Z9b30JXG
DgYLxLui1hkfLUsK7CWirHgthn8h/OtZpza+IhA+UaIgiiYPzQtXoiAaX6KdghfoQs0e3HwBy8xy
UHDOEIE4kWt6NtxMvta9IggzVQ4eUyXouZZjJy45G68GB87zYGCnI083pJHyiwq1OvdBXnuOhn46
buRxLmdRWAjxclkWYDB2eQwLVtVS82Oa2djLUA5fxDX9MR4+lllq7RYHJ1SHV1iYv0hXiXROlKrp
JQTxkZ/b58a6zjV8suiMW5gfDR3nFtjsk7bAgTqFAnOnj1XyNTWyOp1ZJvW5h5l0tMImQDpqaXJP
wxnpN0xVSjRITp5GNvVvP7o0PfC6DtlaLRFUNsCObOYMCo5sWRAUOoyvMXq+Hf0IGymS9KpV65Sz
avp5xP64+D903V4FE8yEj4gUxU2OO1QzT5+CQhcHGBlIXXFe6Y0hf4ty4UPa74WB5MxKD3Jjwp5u
YpSf1nNl9mOi2qh06MFy5TZ7vWDn+EeRDFYz/M6Lc3AUFkHDeAZagUEeydkSm6U7zsBOWp5MCXS4
f7DktXuwfVhZYhCjqLgyz6QaGo2WD/HgNKq+OqHey8SrRVjdLT44AE/fDJ+P0HWBbSIWdlznih1s
S7xd8kn31aD0lU9wSewihdTO5/19j1rG8TlAy5TQRinK/DNsLsxidnGKAJ0A6fybbj9if+4WB9t4
VnMiqAnSrbMzdZQN8YBqKJFQnqrr9IoB+RV6b0GYAAeQ6ueNgzFzSPefCxm9IV7uuUzbt7+0U2If
iVHr+/uVnmC8Vasre41HP+R5KeT3tFVle1Z5LfdMH/gOiNjBJIVl0wU4jdM+kAxbm5pSN26LSLNY
ZqAHDpzyIVhEUxP1vAMiCTmejMyH44XDqwEWOSdFkMAygxlvZjjbRYALRut2UxjiGZRldzG13sdL
k80IjI0sXPMtNkhZyrGYhodwweYN5h7h+ssGkm7C3IlWuX4xMrkJIcb9r5LFrSjsVPEspANzXxK3
SBcVBuiMoriKX0DqjxxtQtZNu5ZtG/DYT/vY/ZIONEFwhq15R+UDfhkvQ3HYpiOTBGpZdG4YtbZD
ztXNQvaLGQLY9uOZMYFjj1TOv1xs9kxnJuqpKj8A4fW0j5kvWSxZf++G8/54M0qR8uw4rQze56OL
0xcOLLyWDN7l+gsQKM4rQRLDe/w2aAcBsIwB6/3Yu3evYvOwy0cK602RmMqi1nYFExxz/PoV5QGm
BEIC2sCM8eqf46Eu6K8FhnpDMi+A4xVlcAJC3OpDbpRDQgVfGuCsp2pKslk4o84U/sCty974v1OO
Cs6rva0/DqYl70r34Oif1e2E47btoWhV78blbVnlLfUkY6TflBbChm1OlyOz0EdvmnBeJii38lKK
nEnqvHItZnAWu+K30oVnrND9ai/CwWBqCAV/uxO0Gv+aS+f8ZTB5z84OewMz1RuVjNalo0w19FPn
YaHe0tGKb/SlSCDGtuQG/4W7mgc3EQiD1JQFdyBmb9MIGyQ+ZLIEYVjXZBOXUQAT2LMMTWJn9bQd
rL/pnHk71G9EGfYrtc+6WexA470Tz0e8E2drxaQt4bEs7J2nVXHMSi1Zzcm1TBrpWABvAulYCgsX
lMRM2GckeYjwcbs8hoUwTnW0vOv/yLJ5A1JDXr2ugowXRc+uAI5G1XYkaZTLlmyMcKpXsqOQM15c
j5vlqdagQ416UmIssp2sPhCjAb4IEVo/yXeKVXcF81qqe8in/duQ/0dQujDt99HMhy04mm0XM+MS
DVHY7acx36ujDOsPitO3dJsS9KnteC1XBNesAN8fhLvSyuTlCqTAAv+Ko9lgR4HddaC2+llA/jCE
zUJuSFmxdqJgVDZrXNOZoDzXw7kRBLFc424NOPc+zZ0hHo1RZ5Pvo87JH3xocaVi1PF+cHcN7GRg
SCioUm5cThwEKODw0auFCN5Y97Kb9WpgQhV0QcRaFIcieSS7VkVXD1qrL3pq8fJ9VoQ5Za4xYh9d
99nI1+b2OJTaYGLqq29lNw59xTf7or49VfmkanBPEBq4nJxB0IdRSqRoSlTv+GAeG6Mmm3iKQWfB
gC/6pxeIAejesWvEfjz6FklK3EhBxHlitMdg9T5L7HC4doZPSODyzN3LbAu+zL5SgP1+C5tSMzIY
3gAgO8PyjhwkNQWiA8Unso7LAATkLxYLCQ19Q9NwLUL1Y3G6dv3GYtjYJ0L5GXTCWsiWJycrNd/6
t+6mEj0/LhNMA1bv1Mia3RmNSSP/XsI/3oU8Z8vv/VW4kp3JprjgWn1xVB/mP4Soogh14hxBw0rs
AcEbbKCHi/lR5/R68nuJfbInnNeDK2qXa8zIdLLH04Z6x/ffPHNUSp5e/rcmJVSQt+MQ7ctWnT2r
DbfnRkfmudpZzXbcdJ2vpo/2nQaeRbrmfMddUAhLXI0QgKuorK56bHboyrBTsdhTfYbuHaf5JNQ2
V6GXnIUGfQ9dXWpYRNsPOExhKrbYujdOVCjqHhUSbyu2uivDcJgDmqVmRxbgRRqUUuU4b077G1Pg
soN73IclZgmhtZZ/BEtD+UuuhaWUY1TTVYbDqmtgyy3LUVO62NvBakigmR2IWJ/SQ9h0uwtsh5/9
ITA467VmtSuDCrIxalHlSnhNs6bq3LSBEOJM6yY6U4W/DqBNLAyHV17GEL9IiTTwU6R6fdyKvAVc
h2dtUPSsry2In94LBQHE1L4P61D1j2pvn8uT3r7dwiZ6ocWTkLMr1X4MFr3l9tErKUPzwT4RnvMM
qkieXhKyAcOfcr0zhWhMdaCMeaONX6kg3Kgb15AzwmscQBppPRuUd5Ly9l70PTgGzgI42/rb+CU7
zRPOwRs0S0aYJz68SiVDEOvDqifxoMXxVn3ojHjC9YMknZbv9AnMFPYkrywtdtNiW+mDrW7rg1r9
ziwXDNJIbdf2LcufNwxAcOmsk7GJUgS3W8iR1Cd6/wZDSR5wIZYecyiJB4xoRIN4XMuJ3mp/RrKB
DONcwkgWw33OIIMfSHMPHzwL/JMOKvQFJeReSx1oQUkxKhw+uqS5Y2m4enc/0NaV420lidDFZ7/1
ANooaYJlTt1EV37xyX4HfvKp26qWj0bIiT/4Pzf1+BlJB92KmaoTP7e/FJkB7aMwvEjxqnlfV7el
8mwhPFLidc/NG/uCJ7ZQlu06dD4hzNHkS8yy2MINdlSHupU4+rBqVwrJI2hzT2mLoUmDbPbAqUw2
YjtuFotIecYeCKptcwhZ4FwAC06CP9MIHcDve3yYfEuIv2hxWRf0xlyTt5WONJZYqw8E+aBu2WeE
UgLjHw2Wh/sure1r2dg0FND4PVdWdwoU1lxId8FCmE+VYWDGJTlC4pulAiQNWwvQjWYKziK3zGgp
SI4/Ap1dbBLInCWoUtbxP1eazrD82SazE5oK88cyfaAXcCDzYFFxVy3ytpR7abjC79bp8A03K+LC
ObPNVQm+XSlY386YmJEsfS7ub274GL04TwvqJlDOizzwOtYdk055Nelyxqm0C5nJDc9r9FzM0kVt
9X1D3GDR0DPjCH0B5EiBh28LLjCc5keyIipJd2bxWZPAn8kpJUXaXkzM/57LajubYTaPkYuqEkGM
uRDtwJOClVnLsXl/iH2Zsg8bZFlbTSDXvmhbpgqDot1I+Su6dTbpfZmg6kDlAss4/RWmFEcTxK/G
xzGMUnN/OiFHUohEaUwQvuMLsNoWDyovze7bOX68ziDSDg8cWl4ZY/6sWjkxbP1fes8vgXk7+5ln
6lNYbHZ+JcTX24CL4PTgw5EpzA/GoJv9nF6WbicEBXN3cL8JBBrYKmgN/rjHy8xqJbSC3AbRaqxx
DOAMFuidOWOazs8ustmWs2vM9x1dt33t/69y8jvK9LOpNZPi6hUGWGIKOeXcNt4voeA4ewT3Ff5J
oAOsBgV/2vM3zQXqdimVYNnfb9ggTbl4eocwiOINAprf2VYa/6Bo55d5d2RfxyDbk3fDr9sVxAaG
dgbdTv9SB3mlqFnAMngA9e8mGycoLwW5BzhHuQK7O7W6uP1ewX7jaIbU/dflhXoGiOO1RofZu/B3
89SwsVZCG6QtTVfmvPOKukvNvfJmI699arX55jwDsbtKrddfFzlkMVWwK0WtU9cAnPdL/bGEzEkL
RZ8rm5z1xgKRF/9svUfpPY2LfiWbuM+Z7j5nf1r4X7WQv9tUCqlP3r1CvrZgwt6wGX14ghbzytXO
TOrC9gUwXU6nLgZyfi1BDv1DtiTPWv3+LH4xOun4RQr3VR1/kMw7sa01nkGCpngcpszY9wY4bcN3
fbfMnzHJl4yO8LhSN4q7FIX/fdxrPAW7taydyoMBdsusDhNPYR5sKuU+MECqrqNBSYWtzrY22oZ4
bffXVizyr8Ha3shg2CSc22whDSJI+aQG6AULfAVk0x8IHEe0ShP8umGt0kkq326Fo14JKVisyP6T
tReM/IYpwmG6erY5nNQR3Em5APE8KXIT+zY8FqnGxhT8tnDO6kbU6XNSjuVu+FEI9mF+h2bakb3g
bcLcPnhHdCmDpgGRdu+eu6WUJH5U+xTzh/Nj2vUv5VWkuT0wewFrARtMpsLuo/o9oS4tO1emrqtX
wHSkyJaUV8laEtVxBKHqnV8naV7iD9eMeQMmR4wIFGgKsvC61nv2IXX0n9iY0wtMs29P5dt35Tg/
7HP4Y/bi3oIv/zNkR3jiUp1rgbs3pSeWSP45ggYWBMCo2sDJaTENj3rs3xZM5WMsrh6/ENrof9b+
0xNpTHn1n/DLBdq19Uz6mZqFB+QILRYkKL7SKJ9mXghp+Nl7PmsTgJY4WPa2lZ7wC3FUPSRLp0IL
ddkK3txuoBovbTIZ0u57ecGJVQ4EDWuwkkY/zubu3hE2fpHabZDFrmbQu6Gs5OXNjFgjyaxJMoyn
nvNQXgB2K5xHLkuagvlJP7Il8V8pi+u3zzsEZEvnSA4mf7Yk68+mfwHUbp8SnoZO+BJbPpZiD3VP
VZupNIuihazNZv+wVdjEi1xsRD8wL+lNI+bIEtiwJt5FDvvR3/nnrufZ0NFexeprHruAqIV7rNc5
qWNFB5tR8wFJTrtOZTht6VDqmYmMinMEmSTu3AEo1vR4uAVWTKJ0U/CLMzf+NLwktaLWK1kExkKX
8Nes1nX9XJTZOqFRzr7PAi8JTLmu7joRqM1IziFpAwVtLc0uV2t042rxou6wUVdyodgAsZ3vVTgh
vLFUaefI7taaMprZJ0s+2GuvbQDUE9cQTt6teZOCWFnJIEkryrrCMPRYoE26sLhBSGapTDBk6peO
UXoAoUa55TZWTx3LqWGvxtw19AgorDyg6nF+t5iHfAyUKKIzRiWcCC+SR9MYpILANLQMwMJJ/pWk
yhtntjcqQfu6wf52BB8wM02EPHc7b3CjLlOUk9j0BIF4ZyOhZ9zvktyopMVRZo5VHGOuX6FHWT4H
dUQlBViCjeRy5KEL1rrQrHTgnlGazm19pVrcp78eC+2uK0L2EMehkG0dagmgiWrmlS80l86a/4XO
UaB5pf6jKmjH15xknRIQor6L4pNValboYqrTk+xJdj1cyr2T2DJqU6PacwQQEFGx3nmTrsIvle3s
Y/QiRmQBfhnkbmrhHtyhUCav63mrzLEP9baYVsrfGrefOkT1mfaeB/aZjKsXrQu8lu8GxFaQbqrT
M6oZ8T3d3haqpZThyKAs4PLT7dcZ+1I6U7aSDeANBlTZ/J9kHg3DD0HaRMvfp+J7Kkkivr2rAywK
8oeRr80kOrGTbWgG6auNQSw3ToecpTjiKrkeeGLUxkx2tbSws/kFIRi3/jbh+bE//MAJ9tf3NZ9x
S4kts4VySkZFmBlXVfnPyK9eKgV4BWM93MCE4s3KiZRi4Nc/0SuhxvfKlRjaJA4FbV8JErKsdX7e
SuRsbXiHAXpBZX80qGig/GHxZLViS1fE7UeIKLuntobaX/1OQCTvMSAaF/qUrT/ZEtcUGUKCkCWI
ZiCn5E2SzmFgJENxprQyjMPPt51wx8Qz+ICdLGpy79MmGqxMT4n/F8BX3hWOT4KUbXasKzREuINL
gTcF2grbga1CVh9dRoevPwOmO8gFU0ZUO5e8uPgcDP354tujVSOVDMXJz+qsZZTQx+lan1L7p9X2
1DB0n1hdn612govDb7xuVEDDXeprJ1x4joEvIsBLDJjc03oWjQUl1AyU7AfvtpKamb1smjiDFP0C
/z2qMwUi5AOW3AW2QAYiUlfgPPHkjOK9KhjNMQN9wNMUm2ZWGt534+ykN97iyktaPxc5KVNLVH8s
gwyj+tPxBSCz/hVAH0jfsG4U4EnYopsQ16NAcIHeFWCneu/kG82fm/Q9EzbfsWmR+CEh4VuiyIot
dUICRPQp8LcAQ/iM54KW55q6IJdpvDy2YOXLFVJVuFEi2PO0nuTEZTHVF1ul6bZDD4SxSkJyuuHa
RuKS5DudqhiMcECOI5I+37jI+JuGS3RGfIBtpwkmLK5oy2uhFqP54YlTWXKjVULpdAUhj5SdWWsj
mKenuYFFPfHVZ4Mej4IYVQJMnQzKNIdmGXWsQqgRcPAlW532auY1ohCYL9YvcxyROLIErj9xbF0D
15C23okZy0G5ATik8URcabUB9kqniasDXVC8j96/qKCZWNXX2pyd0cECgMvrGB5Bxm7UxSZSvKso
uoeo73Yreh4FQGOuoHVQOdz4EcpQ0xQMsutH3j4woAjF60DnvavIh9nFJh3ewfR7B8huHNVS7sjq
MMo6NIu7v1valqzRYZrzS5AKmenHXQ7C16x84GQnIt/cZp2nAkdmPzb78Kgtz1z/c4PCe6ULLgjL
SFKC3bNl2DyGL66SIHAPKS9Mk2sIJydLplS3U/Nb7pCJmD8EK1u+k5l7CyztuN0BqPsM4Sw2izJG
3+3ISU5/NuKi+O8n1ss6sHql/o1TK0eDnigvp+ELrFS33Chil3dgdtOcJOPHV9HU5huX7lQstRbm
FEJ30A456WpEGKjZLm8bX0DAqrprkkKw6zTqWjh1Y04mZsWONo1LQc3EE1DqEMYBKKnymKyvg/tv
MtBGMjJT7Bf9J74UaSDd4hyCu8UU5qKDnYyoUcbeWf0jRBrT0+ihlUydeNPaVqGi7EUr4MVOw3IE
ttJUZPVr0SIHm0ZCLIgwB4uvPbD5tdJ/H4ZisNvG/vTZw5NwhCm20XWRtjKceOaSYxiqEMh4E0j9
5N+m8jfWK67LTS+Wt9TjefjTlTozNQscpb5sK6CkJNOI4E/3Eb6/H8MAfFiG9zKpd9/7GGgwx5MU
UNQh04/Dc0fCMCgbRE61t5pWN/2d2vN5muiMrneGDdNGKeYjVt7+Z5rjMIOFuvdjmWPQceMVKHUQ
CYIZQu3gp/WkKFBpbjHPGVdwXkT30S4KB9Qnse3Owt8Gd2LQaTeilQx8j8j+h571u0EB3+q0Ktn8
vlyG3/2SwGQXGX8wxSeYLZaZk6PKdZq536X49KCLj766vA0fv6s5+OC3kMFxEb4b+/LknTcU4il7
fjcAPNW12qXS7m4XWE60v+7prvvjN9V7gKLaBuJyvfInXkLSGboNHHHAl+AykIMX0VALzoTYwSko
F4QHr/yalA888m3jsoSKNW+ZFllxLWqWu5JqMg//EVP+HITldCdGSd3qVkCMmtNSKxubV0DAhhmI
e9bEYRJ5uFH6g7kGSaG5Uaebxq+Zm2Gs3uDm4MaqXee9JS7qG8d05hyzLZ6tg3Er0s4tcJVvJSR4
a8tSoaYDhQ3jwDpxOzZrQ7F1dGtVVekLJTZrbTDy6EQiAB1N1ISs+lQLhN/vXIc/o1/6znj01Jmj
Um3pS5IVQMhU8mSZ0B3yWvRrSM5/uzHiPEEqYtJ0d41efME1U+1CBC0+NvZvf/SGfjOPNpVdj50K
FESgSdtpAxBJTiFZ/JYYgwA6jULIR7I0Ehouzmz9D903nsCqJuwOphEk/JI8U7eRiUHATxcRskqh
5WqXv9bdHPHzvJ5R+ZZXCPsoYPg9ZL2Vjj6/8f5d95ELzj8GTJUEqu4JJZzbLNEWRh39c1EltwKM
fJac1jhNFKu8ncahrly3A+oPajkfQ5lZYWesMr1qpxSRGRNBr4y34JI92bKuRJpnYwz6XGmZ6zS1
kJsNpzexzQTwwhI8oeGeoECrdAFxmBPJDudbpiisPHpe876wPpLldlhrsykX6uavM7DndzS0k1hK
5osGKqdKYTc6xEdKKKjN7Zwy3Qb6zNEeYCOYVpuoWi0o3JBYyI/N/8UiOzeKio2lyVbvo2oFU3rW
m+bg31oQWsXfsl+3O8QLSjL5d9xIrxzaNrVcAnpsCeaeAetx0avxrGx/1ygf4c2tnLakMzPXVsOa
cds68ckA426QzrWdmYd75DcO8bLDCkZyDOiNqQfhxw4nlKjPDAehQewnZxi2PG/n9DUcQPviTrDr
/huKDVxyOJwHon4jvWXEnvNohpAwtqoFeOv+oE656VXKPjUxIuTvv8SrATBK9dgWuNuSZ1axdx2l
l7ih+7kSg+EPpSMsAZyQB1UAByfLt4EhqIbPb0ovZisOCAl2g/VpXtSd98mFKy2HV5GuJpUuLPJc
4fVC+YpfjguqIUnhgUT3PjQ+fffP1zohFDarljpGpTNbS45I2mfMvp9wn3GKs0hpLZmWXodFAfhZ
ZSLQklmcxKbSuBmhxSzLOyo3/QERKnjJJAj/NuchDtRqSUguhF91ji9e6OxpQhI2sOY6bvzrVGqV
m1LhCHw7836KijvHAg97aZhYfNrvmfq7j5Cp8reSpVvdVaVO+NJgXyCyim9pxn0OTCGGHRkxIpKc
gMzwVaKDzfhRfkYnqXzxtx2otiaNyxmEitZy11GXiwgRXEEik/97tM6kRuLou5140lC/REFa/S17
Bs8mfjIgneUFntbEXmjl/g4diR6RTObHTYHz9fByaCf8sWFrSOOXWvIFXzsVsCzrsA1V4TTrURkw
1yF7znsYklrpInO5hMDpwkmZjMHMxcwvLuDpi2G4gxHkztwiM8/DW7wYq3DLT8tiHbvYSKeNGQ61
T/UkvpO0bvEs/HgU+lxYXLkrUquUuN7glmH/HzTjdhI7bKOH7I3zPY//qXaL0sQtup2UUyuotFis
9QUgULSOgi9aur5babaA8IQqzGOzS6FsMbXNx1oBkNY1PVsJEVvgbg1kOOokf0TxAMEOgFMvFw0P
rIh2dwLXjUoDEM8pzB+Ycu2pPHW/8imLqmF9XrrQpslrQqziJKTxaS/46O8kqUZTokaYz6hm7Bbt
LIrICc3iQvrrPHmvdGugsbCYJWWsJ/adOQwmw6Qlx3jYjWXsjpB2R/7byW+o1ECxCv3p+QVPd9qN
ggw0DC9R1R0cpMZ7dxNP/0UF+9MzoeVGojHUh92lhxm/6Y1kzGnQzCEHEfKnBRIMAup00Wravf2m
FXBj+eQMn1C0Dmou0cWDifIvsap3eKIM01DqVLMMADIxSnvVSc6pyp1m14H2zu5mguQVN6R41kFo
wkUdd1BmQVtxxPnzrVlDgNHl4Trxgk/XUVH0jE6kyZanLpSmNqK7VxLCQyLasZMDn5CPBX2q0dIq
3nC/4x+fqw4ph2krwiB+nkUGIYHl0tqFF1mU59l+KKDyKcXuLybgTIiCzX9Uu4PxxrMFXHKET6hl
WJed6kzaL7fYXN4BAplVAP42zHBHRYayF3JQsT1Kt4GE441YOnZF/0e/9HyvJgk4384OThlD4oFQ
8U9zOAQdGAPrzF75vu53naKrX7W5HCXuBgYdV8A3Duada1fUjPPSkbbATGpfcEkZ7G3E/ya2IbuK
ofokJFajpfCnlgm4/C7wyqMmAVLk9jxuVsAZHNeeIwAKAunZRXDqnYVM6PlgEhrEcSs+oN04Mdcv
9xNzpkiwNMjchXkR95K7X9YJNOZxLLCcPZT/bCxg+99anjpMSe2DSj7+zls8x46vEap60KkYR50M
MX8s1J0Uem0yLScI5WV0C4aoxI4zajvjd3OWBG0cVM+rdEoXmZKVYSMlOk3iKX+ag84T4bjaNjdM
6DqfN8++2f15iIwaxNG1dz1j2oEtf+Vf0C2RqhwxIr1N+5C9Om4mIZpcON/RuHOzgWrJJvur1vNO
Wsab9h33lTZQlUKBgR42xJz0lWlWyqBCs5T4RCIj3f5+Gq5MqYA3ArMteGdUWx4xHl1ntB0Z+N1g
PEW8A5z3mFKLvZE8TpY4191DNh58OzxyddjT1bA6dRjPodN4lDR4lgqukS1ImiIwHSCzq+jMFYrk
rjW6GLySIYqsLTn40ku768GVKqAyGQ/D95nGj/Q4f0SJrML6SrwFxp2ayhrCv928oPN/tnv68//a
u9l5sHrAUTG452jgQRLgL5gKOmYQrwWROj8x/rfnnlvan7+tfFcWkaCDYd2O9f3Inb4gDK+ILE7x
TmfDAUgs8k5t0X202AC+NRV/xrFUSMrWLqLPGkJADC0QbmMK6/Nn8Oy3uncsR6gePU2lb9E0ucXB
gXpdRdLMfj0wF0bbLmKdqWDyMcgO8ycBroQkvMZ4Spy1Xf6j2DrY1LJnUMJsw2dOJFsnLtQp73MT
uNCa6ns7Ux0UUILZqGeA3VWHIkPDfzp3AqvEOusz/JrnXx+xu5+92mE0BnwGGuvLflCQ4dehh4Eo
vVO/D/Nbe3JirBmrZKm1SpvpLjW9LaknzhShhjt7eBZ/QrVF6+zGL3A10YWq4/U44Df03LxbqqtQ
VOiHj694tHyEMLyBu1wxUKfnGHN80Rb6o/LsMVJJ7Uqy0Vv0DIMNKbFtcwfyCkFNndT3MQIkR4rR
T3tPzvBYKyeFODiuIhEZt1TdL3nuUfK2PnCd+rfeb7KYFP3inLDHl18dnn0Mq3tQQuefXXwwGsKU
qte2kN8c0wSKsln8WcZot4alv/sxAIA6QOzQLp6kvzcqq41uf0yGuT/e9Zogq+x8V2YKTxywNvjN
/CMrQ/8glzSPkCak0PjdRgJ6kX1R2wyEVThFWkPsJ4p+6tY2lxInGpm5wuRVfzWZa9bdn7sUH0CX
Gn2gabhC36wcnBXC1MsLhb5wtevSKte55KMueERDlavm4tssGNe3MPTIJQ3Mei5hVSddJwe5/JVh
TgOApAT1UftsJM44foHWYYlX00TInct1qwYfewRsjb5AnaPdSbeaIGuFEQvOc5ZncsWjn3c5wMqy
QUWdLIyD2IPb3Iqp1Mtvw9rsYLcNs0X6dosUYmbnMN/VluD1tmcpzte43qi7fEp4yEghvs+ASQEa
E46QwCGn5nDmhlr6nQqX8wsdey2gdn7xvXYxqbVBWZesJi9Rj8zB8nP5F2REDYivO49BgcoY+6Y6
mAmWz8lGfIYKpz0A0FNH2wluBSzUR9qiYcPVm4AWEKoZ47nPSr2uZFv4zr53pe0njevWjU4dkKZG
H4uG1OffVogcRFLHcmKM30PggMBJql4zg3UvR6efVoMSUL+jRm8awqSfgD2ORe6w4IMgoJJ6fqT8
rlkyk6z+wY82VHUnRn8U4FP4EnHwOykOfy2Dlip02lI8EwDiqjRhGnZdZwWJa9kpw6N5yEd4l0o8
tKUT44ju5v4NWuTGr0Wcq1GpbrFQ0KGoA2wACWxTcuQJgnz46gk2iqviCc4eEOfEw7SjsMMgJdpu
dzucVeyiWXwl8ghP6ujHijXINAzH5BOcy2C/e6Jsy2x+y5hNlG5CRhB+s1sAV7gkePoNsxEgbUWe
dIiFO2E8PqGsWuIJ0UCvZ8ftcPxWFyuREICGo2w1GCkL0jP8G/BNXsY3awIL+UPR/Gn9FGMU72Sq
gJBPAP9IqZd9Oo+MGLHJTKKpk7QgsHY6JrGY1zRw6SLhL/NuoQZiZPokNsjKJDS1HWE1GkqkELF0
0r+O2b6X8NivLgDuFJIDhNNUXbI4nLZMMVhilLFSLqd9T4f0aeRzS/Z15khj7+o8TBHKDPlsL/Ck
Tidf3J2MIUWj7ZRJjPx5peI10+qvjoUVp9sg1+4CmQrOSxwCigXu/t7OFn+PgicAfjX6n5F/ALm1
2kSKTRiJfuBYqO3PlgaSFjQXfeI70JDwBdQDhORCSDBEMLZ8x+IRvyUD6X+pC0558k7Z1NwZ9H0X
yV8yJ4C75zJfv2l4qsvCeqQc1hIbhZs787jPxvU3tW8eMgSgtGjly2OLtOOoQiy48QT1gfTMTnex
DLIaa3YxSCNmMF4GYjM03677sNl9XBP0ck9gAgj0c/ksybIm0Xiq/Ko9WshzrWriDwyLHy0vV2+D
rOuDSDy0E+otVm0mGImi29Wi2WA43FhCnRPckxVHhjiQ+1IL88QkggT4hl7+qZ/z0gqS5HDClyK1
fiDUKzHY442xq9ATCtS08bLs1WyCbHiSznEs29VX5FAoc5UTfM5nZx1ZGuoksE7vZb32qVw1mRj4
2K2k4t0lRhm9hoW9RQgWwqKg7y8t0VSgvx/3BIwS2npa+ZtP94eYpJn4M53Algf7iJNkKTY0gkjB
8m0NA6Fpn57PMym5w1ddo7tkf7ekzmuQO9sDWBw9pmBJX2AcUxYqjsMVLeUpGF+qs3KGhfFb7Svi
wZHJZTiRhIY0P/Ddey4EPS1f5s+T7htmDTixqcnr6w6rbLBzfVGPpR/pVwD29PzaIxu4PW8Txv5H
86JdbIdtPfn/c4bGyIwTjV29VMq4QjKoF3CS+HPXu6TmitZc1XB1BYW8ZPBHbNE9pgUunp7wqgp6
dtPcY/O+xeQ1uTYOcdfeMVG0RPJPOyWfIPl7KPgnErXbWOJvvA55FREg8GilbFiHJfOagdoTCcXZ
tx6XTwUdpyuV7l/U3IO8taiAzfEg4rN8l7NsSadX1uhRkKaqL+oy5/mejMYtPcTH58bmGQVU4qZV
6Dvxp4AODbneWQvOBv+5BGvBTNw1iT63HBK/nDAA6SOXt4EWX57pG/Pyw3xKP3N2+xEfaFfh8VOG
MlmfF/tvoFwvQK2asCR5hbPRIVHOPNax9ZX771w8iiB/diPyZwoF9ojpRsVHiquQ6DfxSwXaBMC+
Q1b2gGjL4M2Y2OKWIxwz4N+rf5++B/NAJZvNM3Lcd1MkJBOi/9oWNZbKm4jX+YhDKUexIRqG/1+d
D5++O3gCsTDc2mPLh63kn39M0RyK7KTROQdBASuc+xyONFdk87vtb3oWNObbptdQ8GpPEdaqOnfl
HXwB6Qu8/r4E1BWYmhfqsxWwib8BxeWhTEUR8194QfHtMY4+YbPIm9OEkF6qyJuqu9xTvYNfKsAz
aebF88ATesZ6ajWMFmqz2R4DlrPLoT6I7wFlkrBuM4j4UVrrOhknC+SzTtnKlgOXB7iqyUK4NaEK
ltPrKUyhJ8Y7eg7kUtLLazwAmANG7eTX0VD5AkkMZWovVhkiNfvKOb30iT95bsto2tp5FekOEYYh
JTf/CWmlMWyuSGRl0MSHFddfIHLA50FBBOi5Um6Rwu7HBHnA8iL6l9JJ+L53iBqxtFUtHYTe7lCW
UXS9Nohsf4yihOi4hK5Lw7w4kdRqFvviMw8cCOqsRtu65PEE3w3gZuRwLZTqZdTroQr3e5+Qdcq1
B4Sr81iSuaeiqRFbEpKLnYeJCFQeW8Tj4+exQ238EnnhjQu1SCaItTz1b1dD4XIjyqrIU2SZ1ynk
Iz2agMzfNsbacUOK6lIRkHxsCGeUBKxRIVknqw4YCT3SGDDflRSpIzoO1xrKh59x7CauCSvKIMty
jAEMxrJvVJOxEza+i43yBXQP/Bn4SH9r0aRUMkaC6v57I7KJ53jOOJk/gI3tfWjRWu/MuAlsYIsl
kjjCbuZdnqOe3xBmJgsxGiDv6NWkHYhoR8zA+3rmy2msZDOtsDwruMljzGkzkIUB5npcwaf3AcyE
MiKL9WpYVqodQk0ULB3rw8Qgs6np5LzcfGG+iLIVa+VOTxWHyeF1KqydFQV62VOOPFvL/5Gqa44E
kJhhNgpCqsGhUk9xn3lMSL4GKE2chQaAc+LEAwd6zPD3+j/6V8F4Djj/3gGVBFZBpGy9eoV7wC9P
7ZmijEtgJDwrxxPFu2x88jXj+TgbBugE9vw/I+XdMtVOxjj8WwK5aRzbAaLn3sHYmoBQO8N0H1Wq
ZDbUHc6lv+Y9h67jUGUBVOYHg/rrHRlK85Ut9FCKquR6b9yL9D7oQWu9QPiTvpHseoc4Ft6WViZT
WVFcr+d4kqWH+H1gjo2DLJWklQx2o6GI5pTW9bGhdFUXYKluIft1fpD21eFBBOSZ1+y6DQjVOIlx
g/9iUKSisk5UCp6L+pgWrZRdBsdfQNBPfPrjLUU+fMTX5aXAPgikOSTnLlK30Li2KO3cgq6tpe4d
pJ4tliN+yoOmwt7CuDO27ek2KrJV3k5W09szCqdkfzmIxFj9P9zBU/U5MLmo2P8YTTdcvJemuTCY
xmsl+vgxhkvia/hAK7uj/QxCm5te5JzpG8iXdRJmD6+67rZsVLwC8hjhYcoWSI90GvOPICvS66t0
GGnMKRbcs5K4/N2OI8z+vBNwvZyp0FionhBdRt0cqJK7nZ2XGPQlSlHYbfv0/R6yVFOMJFSZT10c
e9gCGB55GVaeWIoRXwic61C6UmfbwsoyZsx2kyratCA1Ao5hoUjPsOmC0ASaChVlvQVmAVRBDsrb
BtdGTLubuTyE3vH2jbNRGesO/6fFIM8ej2dSWhZ8OLTza9B2za2cfFMjc1E3Wo+I3doCol9NEpnS
JoZcVmNeosdYhWZVpt/hPo4iQY+B72Yjr8r1kHwp9aQ7nHGe0rbhY5KMAJ/tHjNvl4W8jwoAJz4W
dLa7tl+3U2Sn8J0DcNh0sMUWg6yFOLBkQR/a6kotEon4K2nVOnhcQ8V9c+3cPSrxGcsQ9F+tZ/Z7
sRU3YgLBTjDn96QlHw8jKt0Xlvgmqqi8ya2ujmfRkBYo2W8XW+1Etww9fWK3n54NPnTz5gviVe79
qvU70NPVE1qxFwV+63iMXZwP6sJSBL5S4c5JGHs3NeWGhpjnPQQF7dulT8nwqTzeXpgNbAo3oYwo
o3URQuAyvIASB7TEsRClz5He9m9McOHd2lFvrHzAnyaj4M6V4zlInF7mzLXYvOEfwcDqCWRQ/gf7
YkL2TUB/bsEsPFeblir9Aaxkd2Uy/WwcsBBooQXrMAZv2F2MSntLwRy+goN6vLv+vUAqv6nykxoD
/Aya0O3PdT8c/b33QIXEgRq5MoSM/f9U3uHzBTMgpPzhfFIJ7tiNKNaSM/mA1RPhPOKqUYLoj992
ngw3dSXrpdhdw6lQHcbPAcPfMf7g1lS9h4daoDS3dExQXGW92EPTTrZgIL8RPW3EU62nJC37+wWV
uUWZXWN1kxw490jlE10RYrdQS5MY926vA2lq5jqGAlgWhqri9gWo7H/VAC6T3pkblQsZ+NsjHaCo
6Sq2REYrjsTudknPGTRevJvSQgx7Hnlvv8ZrubVswUnCu4wMDGd5Q+ajFGju2NZ0N3GPO3ZpYh0j
XUwADSW+ovhuJBRv9IpiASiq4FlRyau696iJ72xp+GnqlJkAA24i1okqB1InKVbKJo7nrP2lHWEc
ImXWrHiQ15qaOP7t0ZWqFygClTM6JlPL4NUo3NOOmxtGL66fk6OkrPmaXYQfeT///acik24Fy6Gh
e/lC3qmTmq8IiY48j1HVH6vrFEnrrkWItt/WHo7EgP3AvAz+lSBf0HCjsYyvL5B0lAUwHw84Nehz
LgXNn7dYQ8kFX9B8snd1XcgRMBqEbZkKsGhr8AQ9rWfCtXtn+JwyPJtxEWpvHhXAlT7P/Xf5+1gx
jQTuRkvEMUFvjUDiJ9izOexK77KAIEBXWtwGopGRLW7esBy2oBqBVEhKhv56ngM0ZE6vHSgYpM2X
N9ADkS2VElY3axnbZd80Mu4GLs47tmjywMftaILXM9u3+lisXDiCdt96uSkaXmsI6IsfXepujH1X
xNL4y+/rrRAyJ++eWKGo2+r5fSe9q/I+7oCVLAzU83dvVqHAh0qxX23BHiHCh9/1Mb8Vl9KrT0mn
FxOe9MVnphU5BHtAFOSSLzxOqchMNgM+BtbCP387hQNkxaOGRa/g+x3tpsSKDSPyHnduZxDZEirh
IBh/dY2fqIaNuuImHxZsl+F31YDCu0OYs4X9kRy82sRMNcsxBBaryafHe7SZrwXCLtKlK56on0S8
0BwrOLSylV1Np/EZFdcbcfAD3spKAh3uRjk33X+K7Is7IQps4+9oGRTS8/NTrcoi5tH90QiAwc6v
q74yrtDDDr0+SOaN1VXCoyURVOsFl2+8kdtSHb/y96K7Ws7N4sdIbeKx2Mg1OcvlKia0/X7ictNL
qpIHmPiuQqyixy9Ge7dz8MsDpnlRrdYO0uGMDLrm0EMSIFBekDj/riF80+Zk2Pzakg97jHJScUWr
rXNj/gMaZyUg+FEF+3TBr64/MRac/83In3rcQtaqsFNwX+fnfw8xxs3DBN6tk0J56Bb28+Y33UTs
WyGbHopelRRE7tf+gOTzKHGcf8yxlcfr65EBs5TOO7E4AGVXlITrOjD4mGimaHJQzzUcPtrX3O7r
q6XU3rFgrYZtsp40liTZ43EbedR6a5S5sOFKH1ci8LhQ2GAo6ajMfQ4o+sbiSQkBfQo0tl+FZqsM
XOaBAoS6sl5Y6FqnLHXDZdprsomgVVxVl3wzaaloGBUcBvqn/F2T3RQW/bcoaZdSQQmorP0/vhVf
622g8vJ7XV/55bwN7dSP1j8t++4c1nDy9AbjN+SGoA6BOunJe8wuoY8XboyO6q0+DP8QR6ygmB94
z8CRiwBcFKEZ/97hlv9GMn2Zi267gH94VcKTuiD9dGZk2qlkNk3FjEf5CfyN1G8+/aK0GOOcNVK6
TcBXs1XajbQAS4wVyuz7CAGqOO+5iPM+fIYE2TPTLS/howUB/dpgV35MIvNXaen1AZnkuHBVIUtn
RvG055IdEYS+EZlvQ2FxiOVDpOHdoCpLjotcL4H5kTZVm0RK8kQ7Y9Q0Xyva3KpOfr+hB4E57ecs
cpEAUvWieZlWCX4Dn0/E484iCsOHa8GV6L/Z0J3xOS7NnSJkXh6ZtW88FtZyrk/YgiuGN1zZo0OI
c4MHobgTC1jC0XSZV6RCLIAJ5FRu7QTUtvrzKB+3BRfGqs1tQIhDfmZ4EfPIDjbTaiX81chgPvev
UjF77BtlgPjjUIpasQFfmpR9apd9BQ1w/zondi/G+RfVE4zCldx+XLYrKAmOhiXpE7uio2K/hGdf
oBwQmMuZp7+OkqQvwZk16vhfySPlNoxBhjhp40nS4SRE/y7dm26fG9MREEX8vADw5aEZaI79dSyx
eOIlShNqONAni/ilY521sGlkFw4LxfoB0KIQKvJ0HTemiGG/O4KKbYU/3DKdEIop5gk8VuBhM8Tl
QBL6zC13ae2yx6WTN65/6mj/a7CKWL7c+T9d2IZO+ggPSNXgTampQFijRGiHjg1QBOkS3FsOuXjp
NR6TEMDh+PFyuKaT05yYby7w7ucyX+QeNzXtbxebz2g0BldW+Q7dd8Trle2SUIsig0MwsZUDLclL
Xlu5/Cs2eN1+8D1WajBVgT+9d3L6ssgssTVtM1yIeQi3XQo9lwkyAdKYvekisDeMlbYDhCcuaZBj
cTQDCCyegvkJ+X+WGBgXwcHKti9t1D4ne/3248XaauM/0E7oo9NKsgSMGSRhEhw2ZlZD0ZgB/BUI
brskPMijgCJwT1THnESqmRWgTof3zQevmiD21sDbV5AdSfhLOHTKlSqrzMeKx8t2sEqg0wb0XLCM
jw7h4CVeAS9Dai3S3x4isPlYYKXxOhOATpLnJturxWGHon7nGyza1pfzvj3nCjVKqgcDcMW7c69w
rvCFOlDx4KTWt6FU8Vo2OHmmdXdxWmg8qLSkfTM5Ij1d8T2OKlLeHb9Z7pzbBKZ1UcMUnFjiFA5I
LuedyCLozrPXOVgXdfoGkwon6nQjnr0AIqrsVHbqYk6wd8edKis+nhk1K1qav4lkbqPdzY2zPan9
VUqBCzV0awCAIOg/+DhIf61ynGocZD5HsqQGxebET7OD9yQAPJpojrE38vKfvFnmi5R/xjqgOlz4
JfAngSvKwqcjUAFBpjoo/+o2OT/vZc7fGlUXISurbF/8fVVbVZbIYoW3OjLPcmKVdjdB0LJPG6cl
tQfI4vCjx2jGcEO14JXfHX91wpEwARcFo2yTpdRddzmXHjzxk9GYH2uCiT3XGuVVTbYXGuy6uRA+
ye0ONtJlpiLY1isbuK5KgpCGjuA4bvioETuPqA80zq40R3z21nyDFEvCz2WhJYmf182Engir4g2i
wVJU7KNAXCLRTja54J1x7ZBZbn6dFGMhGgdFFo9tiObno883/C33J86byOFvA+/iMmYs7Gp3ih3k
EidO77f7qkmTjoSf72bb2oq6vKtsxa/+K3y162Z+GqJqAb4T5qyxSxk9OctAA0z5tVru4u1UpZMF
WYS/SOYkAoVbUQDKbwTfOWUEeVUV1ybJx6zU0ss01q2fAg7kOTAmnF8nr3hK11XR42QH8EPra9zu
1Nt9JSVJTm7yNiLFhtpYOAbj3wtkcu+c3BoJzmAWYiiQcLK8OHxExaeA3fiy8p7rRc/WSUO9CEIq
50Sm8FzQmY+O1qHm/ZcoIegVs6NZ7y2AdNXlZKVudUm70LJ+xdRQpDqGt1UfwAvjx0bThIPsF9Ki
idxcsxREWkK9RlTodFw5dPJZouxY6Buwfpfm3VvAB/b8Asw6FoDahYiuvVP7/xxLjEwJZCUCcI2e
jOHKWZwp4PLxBGSiWU1vFnCZk3k6awKfTtwnu9oU7ers0NivKR8VgyukbxQDq4ICpj/IKw5GFN9z
NwSdqZEOJCI5nwQa0YXGlDpZ4vZXvYJB1n/szlbK8jDMEBCE+IICW63vg5RLAuAwr+lBf818oIT6
KAI5tvKgbq39vF3AM4/s/PS9M43055jWwf06OuzVxBdKR4DTHRwkn69sT2pnM+FqU6brFhcUBEtK
79hDqnjh44Z8OwDzGZeuOT4AgU2NfXPyjj8NiEkOAbt5JELDHlOcni2qY9a3rvtmllE2hNT3mjqU
BJop/tWCZ5XCn+0Pj/2y+dCrk8P+ywBlm32mqBGupmcycaMm4yP6maHhj6E7OPyKX1PPeW4pFHJk
onhLXUL0i2x9d9PfF/C78C/phT6u70J0BxCTN47AuGgfjMwh1BHOyI5ks6MEG0UxnxlX4KyG11QU
rlpcJ6C3nsrJXB1EHBTTRQANaWrEWgRkdJqT3OQEgQ1KWCY39lv4qiOy7prgVtKSsNNo5s/wZBYV
anXCjS/neJQn+cpHwtwiumqoyQz0uBaSqG4BBwNr2HrDyMbKUgvuGjSvGxTbJfN89YL3jZoXJVXT
Gd7mG6uxVpyQu6uvQBAat+TdCOsNWi/Y2kq/J3gA9kXO1R3iDE2/ARzYpJ6Z4R22kyh/2vD9WvSl
Psp07UWKje3z1/8/DkGWGjKg7js7Li7lAxsjtSJDkxV60f3vcbH2wqA8nsRUST5Zb7jBALcxq2oe
e0M0aohLrOwAsB8iXoya89EWKSM6iR8XEcGxB3hKw+MwDx1RUrJZOw2AyhAPJHzP/inDjVCNfsXY
rjrkx7X/lCVZn0iH3ePE4lF/nE5Kp+7qjfRbx5h/SJjICZjfBpUzlgtDqm37iDv2tReXnGGrhwjz
NiiqVgx8WS31oyayHRxBLOKdTrJKdH7jHCDXkhDQ47P7uat/dq3vg54I8ggNbadT82MdCdj9crgI
PIYtIWzme2wc8RWaoa7mdgGg3chJIrHtYZyCWcrUVVFu9HCuIQi3PYbNmXnDAZQBbU/wOGmjLiQ+
EuqwPoAxL3sLWXeRAlGNjYVwk3tAbzUzKP+qW9mh4tt3HozI+16zsn9H6W6munLqv0/SAFI7PFcU
jqef3mJNEcr6nIOFdng6AlMQf5RwAvgSM3D0CiOqSvF66LHqJKUCx0LZUpC3GmR6nOFhLHmt6aFc
J6rC8re45rvdFrHJkpVI61BpT1+WCfLIO+mhT3SODPA1H4fRgpIPpKfYmQlqhhoJo7gcy0NMUCz8
ZSEZFw26X3MFmnn5YXZKHyAaU95y+hsSU/ORFvFZwXkjJkXThIw2RZfS4lGmzX/6zVkgOHNrUmRZ
i8BMX1Ihhq8EAzJP0CkHapoN/nlv7tOPrMZfvOXHADWw3wXmt6nZNb6aoNjIPBEUj1ZYy0VhyVwg
YVWTiJe4jIoLcD4kdIdjTwZoULqa57cXL98r5roMS9RDvUfkm5IrD0XsvBeqD0fBAQiKiGQeL3PU
NPQBPo/Ew2Y903DQwVsQQyiF7V0ds4ZJyrrvTG8E+MLOWV3aFmD5J0dETchZUI1XYKJygJT/j/4Q
JTluV/y5/qL5DYfDXHLum2yBY/2yUXjAIjTsVcHMxTOBaEpYLBuEMFOoRyEh0O8bz7siasnADv31
GXe+QCWVTFcpDxAu3VTwHAC+yXyw6CrKxdX9NptVJLrvcKwMScSbYBBaRgfCK/uMIdob8ZxhEgyF
r9mX8SEeB0A6MkTy+ztilFHwkNQC2wEYLmM/+ku/fcZTqPkYaqHK/O6Ky0yCsJB+HLMLE+Nshujo
2deJcEk+1Tw+1ldiediOu+wz0cT55Lf+fFtM/LUhReHxlg9i3AfAuIKoiBD+mJ6BoZE9ylFwImAf
EWYXhsuIHzp50NGV+Bt8ZjlFeEvW1ufkviZD4lUS/xLcohqbi/poQvm0nNLJ+hz8oLJ5Pqa5k87c
R0fHSmrGMW0U8hx7iiKb9b70xTNZwivaBwYNGihd+zZzxFd6mJTXbcr1cEWEjzfJfC4ybWEYT7Mh
Y9G7DSBuw/AXED7+D925Kfag94Hm6GN/BhctOjAWljC1VTP0+VD+vbVTU0WNQ3Og5YpfXg9MX1jS
wz/sBqH+U5PaQhOlnbNPx0IuVPb0bmBRCMRPnlfRDa+PN6BPpsjMu65jGRX3OrMoS3mRQz2QEo3J
+WjRWTiW+5V5ZSkcZ5ZcFSngyuyTBiJ7hzHj/fGyGnPuh1MWC6DOl9bd+eiDpYFv2TVJnElNmbB8
gMSAs+wjYaG4BxrzUZ4ZM8a2MTagTy7GHwj6s7rR39ILZ1qfC98C6bWGviQEWAtkRqlPsLWTarDc
JboGKEwm7HF496GSQLZvItW5e4Q7NoMCnet3uQBluV2k4Z/sO0z3venvCpJ6eEirz7dLla9bTFwY
tPCp3fofO2bwGs9OlnlR2UIe5U9QOMk/jDaAU9CNM9YjVYlPMAi9tld0uSBQxnCeAfvru5GmpSBL
ft4GdxOiIYqvWhBB1woFKijtPCSPIjozy/hSirT8uXSi5NO2hPQ8xW8fO3obHLym44GYSOj0hc+s
eMl1X2FgqsS+6iKBSxFEQHRAvl0maP7RkCDhbS9P5rS+zryjYivtjtVz/PP0H8g+9CKfNFWpnYGv
fTwGHrYHXVHen1cBuwor9H+JMmywna9Fm2V/rgY8veFs3z7ORN8OgZakH2J+oaow3SPCAC/xCR+2
IWsR2N8FgYfLfAycEZgej4QD5KEjKh52kgsqhzPXgCQdrQQA1F+rPJl7l+qhRZKPQ3PL9TQBslwA
aT5gB2UooyvjA11CvSzEWS5G9frmCOqWFPzm9wVMYZumuFHW/dmCJGiNIYAwi8TflaQ/QOklNpB1
ps4TcODdSermH6+DNP91ooqSf2bJtALL+98pEQLX/UGkYLTbRbJj4kzu6pgB04ic4nTHTErzkI6r
tDS9jxbBVw4C3QP9RUl2Npq8zh2bwQC6/QCWgKsaMNJZqApl1Ybj/8Xq6wlqVBjkbKr11OV3hLtX
O8uQGnz6b5jsna10AcKyxOoP0P/L5qvkTPSA4HctxYlQe/AFK8mmp7wKGt94UYF1y7UvUVKIanx8
XbHZC+ZjxK9PSjDn7+HdLhBobVj6OXzTzoheH2l6xGNGJeQV/Fnx9FSf7NiuMJUAL78XR5AFNfZ9
3G6G43W1h8MG9MRkEvoxU1IDnkNuXcx6RHzV51HP/zUbwTKvgAXLJ084kec6MxaTiE3ULNyv5Xen
MVR1VJ+HC5RH0w/YFhXu6AGFgzt/wBYeecoh5TrHb2x8xiaSxQNeZMAiAvDD7z/wZ/HEMJ7DHipP
3vrI/mewmwZ2fiIiyYYfEu/A6/4JkEOWgNYqVBnJlBSSLda1DOAl9XNHX+X5hKimkbezLnyS0fMY
cS7MP1BVtRJdZqDubAELY9U+UVaaff586sXrGFJQ++k+uyzAlqhoPvgRkZRzyARVJdepuK6r/X4n
TjfP+wVxKsn0bUI/9qlJQfNcqo6TxosPMuq63V8w1nlopSkaz846+fghq0XCpifaLkKl8P9Zf/Rd
jMilKAaA+4tcjk7UgUIXBy171LGMDyE+3B+fyzY5Pme14OJrmBiW0wkyP7I+ipcuA0SKXrq5zigx
1ryBL5bcrXM6sVGpAkM9YyFqUki4E1cgOl5fUDtRhwY+fMRyydT57isP9pMVW3geqdi8/3ednhY8
OpxJ4VZ+aYLGmN2vgrelGCOq/S3AUNK80+iofRPMw1oO8pIYu2ytTTYWYbq2rUUc/I08P3qFLvaP
SU+qtfP9+RFk+K00y5sYSSpk6eAQGnaV1EgNgmMVwlDx4pXzLxzpeVe4iYMEWTR/4Oee3HKNFgoD
/a5bW5nab4d+TyUAVP+P4N8Gfcp7aj9gfdnDv+/9SJ81UcBnTcBtdrZEvwVv/ZTSQvreUuOyS3Ny
ipAab7eyZp85CugM8iarJ949enb3UzFQQMW0bUHCkwdVzZFWypVsYs+KRj/jiFWpa+0sT/YFb1FY
z6a4M6LLUsOlHwk1cll2X2Eo29C+l/Axpk/VcUa7i5KDSCuSbZs6g4NR0UA31QVSOFn80c/Kvneu
LLhZMTx9ztloG9JTp+040iDWyerh5lR63BHSDYv8bLv12DZxq+JTpVvuh2cGW5vnqw2dNyeG6NNt
4CnEx5p3pqH7bJIxeCdhgtmVzj+QcfGMQS7p2qSRwxOLN275c0jvoEMD5wPpnh97DNCweYrNSfUz
VCTf8UH4ejZlRLThPt6BJP3Un9cnfoxCY6X0YroJXUqSX5oL/MeiHgQYiBOLGpeoNqqrLNQw+vUC
NLPVSkNKbzwn57hhqsDh1v+oC3eb+28sjJUqxPYzatigLxYnPbdFemQKy7T6z6cOnGRmtM/yDG7S
pgeOpbvoh8DheJh9ZrSwsNSTKRD7IlIzyTSdhkbMjr9XsPLfTIDFAVC2ZLZXc3OzaIFGXiQ38BXj
jrmXKxlIs7HjDaygxoto8USaevRSFPPa0eC21bkrimTMp4Phf/u6EkaAWooJF6A6GB4okV1oitT0
8yEtgaK3F7esaXF72PBa53018u5oEPyaylQlkHp4I+wUAbEhnMmolVI4PbUakarmc7ncdvBObxer
ab5gV1NUMnNKOZpLdMRlZwyeaeKBXCr5UHGgtML+7p6e2TLlNhrUlYLuJrDjfqW4bpHPJXo2nvYa
wi2SPp+D3FW5Y4hI0ua9fzI0TYjM4jUDKyvqgI94WO1TweeP+INMsClg0J4WrIg5wPhnOymDdT5Q
KwGRupg3yHiA3pcaUpRkODIB/LLoOO9PyRh7KIGNUzOCcetJOe2YxDnEH4TE/kbgdTMkVjVZGlnf
O2V7rRPPH4GekQI06WhaPO62jh3j20EueZPxmejef03qkXATEpkb9fArw33dBlY3YkSyNknhVRBW
w6gmkG0yCzm9S2sqZaU1ld4DYx+vdvLrb/7bgNgrLbBrI9207jcZFiWCESchOIeWyMw6eiS24zWD
GYdQU4bTlWAObog+x3cCVkpJxXeuPz5HOkuJ//FheVqCvIYtRZI4w/hrgCIk7jrK/HWwFdUTfoB1
B0kYb2Dmfy4+NPNXXs2JpbWfhUu03mRm8kxgDF0b/lsA/FxDSKvOrNqmZgkubQfisSq5EafBEQCn
P3gbhbjrUnuM780f0HWhlEb0E7mVneCRem9ccdtTC77ygt847TvG9BJ7lUvwEKHlqiu5g68EsWeW
QKQkNtXqYKg3geK0nUq9yI/eey0i+6hys5vXJNv+uVa3JiFy2x7d31kmDN/nxABtrekYmWoU+zZu
tWyifE/cEIcxvbySlLBEHdNLYweZLGJQjV7NqxlI9KZboJxgyBsihiffkuz36JQUMQEJODRqv07i
YXiNUr7TpAGu5c8UvACYAUYKhHKB6jzOzUePuYRBMZ/iBrB+R9xDqt2gDwRVbR/Ow8OvE7ZA/35O
wzRvzt36OaE4IEiSdy0uly8IQVIYKQYEELPzyPuHJ/8/fBI7D20+m314Ta/3Z+tmP07x9KSpYWxr
bXwCbjnw224vcqG0HVZaedJqwrn8YRoXyksHcyYBbJK6misvxARvuHL55Ys4cZ0L+i33kZzEke20
IKPzhGB4ZPGKMTF2TbohNbzXr021IZgc2fPXJpSxvqXnt7pqrz9jt6WoiluC8jMTTbz9++htQ+KA
azMQ0qfccqu5hNP82OxGqs6MJWvlQ53C0OujGaFbGGGMWP8nZDcwauAln6ho+5DaBO0qdCV3nwkU
N3QjEBjo5wdQL3/kppeCJ2gPtaH1DwMcrXmqaiz9b8oJsGyp57kIl7R9Fh1bNRSy5CpXdWm4ODWE
SZAQRRGu7w3/U0myQD6uDndeYRDJapgBstnEofiuV9kWnm5bbJdpo8roG6ammMkV/narA1u4ZCYx
2tO/SUqmCjqc1LIA069HAa0o0ncWR3kDP4sDfLeqLfUxS3ch+QNMI5IjSerYj0+33SAIIABMHeLB
FPT9c1nFuInS7ZQREQqUKM7/kRThHK2JPGETrluG4U/qqwTlBYe6sWQ4DXuChbnFyBtIHUlgugK+
q27c7aSbB/eaRgqNTGKd+Rck5ME1RbGQ3jp5aiF6rV6UJp634gXV68dD2HMROP9wSWgnKOCDtK1y
jjuh64AGFYpvOTdy1x7Ze1b85mZCljXgJCJOF8jbp9T+5g4DVwJegjMCUhoPuGY2xdzuSQxJpFu1
wZE+JZPJKO+xAiuQFOcjyOFlf7yUkoDrSamYwNhVB+0llz8XIP9IMSvCVIkwLC7DSCSnYDk0sjj3
OyYjGWlO74pmSEY6Ve1n/+zsYLPwUdPa0Ll0SxOqOwqTKIFoaR+Vath/cVHvX415V8gnltftvYgM
os+BeCSunvKn667voeWTuFAjBkPaAeoR4vtlhjpM6uTY0BrSsskMquEgurfJJgwyt+7vY/awQZ0c
q/sZzmmZfdQ0XguKIsMUeXcVtCevduNn9yDbNVimg3YMbOv5L/nWapAZArFTkt2tFE7XOyzQ41Vp
eILKxbgrQGpxBSZaNimOBLBihLbVcqkLUbmmfxqvYogaL0FF4Eew/KPXU1y0eH/Zo40ZJ2h8VaL0
pn4zHS7QO7p+nNeb5Ky5toanBIBaR/fy2JTP9xpuAekSlyAOR8ggEwWmmKFVuA1RNmgkn19/kC4A
QMKCATUzoG7L6EnTFz2kuYbFzhktfThkXID2G0ZbrTg++SQ5PHND9fUWRvuzfpCohI1TipfAqzJS
xG5bFttXt7xyGKqS2nxaYqpe+G9fmQGWUtdpohF8F4NnAcGON8FA2HUuB+ABR2I6oWflW38IXL/B
gXmb8dywIfrmgYOBO/nx6L0PavVVLSeZo+tcJqjB0iKaWnAbfyIY0kuBPFNgld9IrYiS7sn2t5/5
bIDDoxkKOSqpj4O6M0O49mQzCOZHXf5Vk+BUy3RYR4dgltABE3nVbSQZ3Zvjy/NvCYLqe8UK+kdY
pZ+HoctTxP6154k1zh4JSf09+LJ5XwFSE5Dui737Mmv8sG7HNTf0B0c4zQ1kYkOUo5s9nf25EYCf
qDoSzbjJGu8XjifOoFMyA+I0nBLz+ykcYF2U+mLKNeGoybaQFwADg8fFPMRfqU1O9WxrE5+ryxIc
CWycsVTyYEHupOjvMOIxWWOr7515PiN/EmFa0XlUxfcjn+A6irV1DBSlD9/83Pdh9GL0L3JsKhX4
UJD0NaU9WGwXLeb68f25qZoqJLfcB0GcYH0lLwek3WO4UAWDU5UZndWUXQyFLXnnxS9bnqKcAn6N
4eJMzFPtBrE3Kxqkrf0xgfPahYyy1Zsl5lz3MmP7R737xw9EKw5JFsX1bGRlPuLrMOxpDnwj5Jul
UZkXi2xVyGUy2hAYu3bTO1l03J/N1au8bKnz1Idf1voG+WVwVJVTQR/lURMY7oI3LwKIbTer7iBo
vxxgLnmYx45mXjiBLxe4QsVvKFSEkyNlc7xb3oQvnwzTkt0NEjIGGAw4bA/w3OxRw1LWrEjsaHyZ
zkgZuNnnys3FudBuKXSIqf8+J9iV1YP/L66zpBOhCVV5lLZebXv+Y+OcIS0wGUPQq62pDqNSBK+W
rmtyFzTaAw6V1IKpYMwrz6JDw53xRCTPt9j6089bUMJSzkokYxjfS8zKXAnILLiIp0UdfGALkhfG
b7SQY51uKK9Y46JNJay3GS0LhBX5TkkT6xMy8gODhDBOx9zTjfg6yiaEdUKRsKvyviCNphHQPGpJ
6FM/LYfu7NKG1KKJN66eCChrOrHOdXt8PiILPOBfLpH8vEZxqaXN89tS/XhYmIgTKz4pZqa6UV5d
3ynoxAKyMImAcp18u1v0d89EWkpzaRo9s7oJM/liX9Qo2UvuewBTeZcv58kjNz+0vGAsBfNMnZhO
mrQ0gHvtz2UpO5Z5zLf/SVvtnn03As4Lm+hFCZNulOhJJQHS7rYAUHiH5qvaqICk2N4+hokAz53g
zv1ST5xJSoqDL4CbUJTlfdk/+Sz+CdJPsLzuCcNysqLS3+ha9XV6cQdOpu7XE3mMh+mRgOfUQEvr
F8tApWNcjxj0OoQa/uc2/6w+Fy3UazbydsTET2us7Y3YsehT8PnUueYJdhYC4c9RT2Nbzzu+F1lR
5+Wq9fS3HIereN5cJVeG9RTwmLwC3LOQyiuyFwOllRzQpz41y3sIJuvUGcz4tQ2vAUErig9xe+aA
zwfcabEkVq0WT948WGi6cO3segFZG2ZZAY0Yd77nYzcyPQn3VlEwWFQfjuE6mgWGEF9a+szo6rQd
hx8WJqZcn7d8ekyd7CQUCgTNc16KF4hv0MytHCCbrbMFdj8vnbRFuqvaC8mUPx+TxNAUhQWPCh+H
JdqFD4fJ0YXDjHJy4RpiQ5Zp348JptNd7hIjX3ixMbjTpYuGCwSlxLcV4IzfQLIf0o2tB7zEP2MQ
aC//mDw503UBC0pLpsXRIqkK1gzIHzlrqWmVS31oxMar0APId90CU7Bb+NpXZ8Sy/LP6iCYvHTPT
+9lQVqyFbgkYhqA6oUjWGHLagxKABU2cPs0NQHSg/m9kyBnuhIm7CBxl0gRCZVJW+JIQxL3hLYvr
4q1a6nQuymShndWkzQz/sBzPQ28QVPMmWjO72PsSWruUKqhU97LmwPgf7xlt6KOpqqlg7QzJh+BX
nxlPiteE4ow38hnP5TJ6WaTJ0pMg6+IJ7O0z8Aot87Sm2Ui437HeqXMR9sjFrmQy1iYT79SvZEMG
CgFSJhTTXpCkNsLdD6fSNXdovLUnw3tNSK3hr0VR97ohbAUHw4hu+YBUa4FqNLluZ4AGs8G67gNq
yAHbc0y0Gz1bVcZQzctIEnwPKVtvDTJ5sNfFjwXzQu2G6Ky5bNzyIPPWsOROYbMQnKebb3w4ryOD
gUY5X3EsX8ngF17FzCrXLn8s+wHmvgE1fJhtXAdiwa7Ove7L3woxzLuf6aLLHbaU0m1EkF2PnhGP
bbGWEhgrEL1ahUZBqxu1J6T/1E4QYNCUwAi2S2purmPkFYuL3A9yo+7YJnQ2P5PisuKRbrTYjPLt
p//xhuWXKxzBbvJcXpfgeyGaOXI89Ykv4gunBR4j1gFGPnAN0jOXmBcjSirO8TG3tmtbfrAILp0z
R+jE2k8/06wg0An5cJegUwfX7d481SkUCbExy7kZvI/rVk0znTiInLZN6bLdTf17VN8Q5m9shYWd
MjbPJAIFYO2qjdIP8K+S8oJioMd69RhCUpAv6YPfhBrQDLQ6nDQHNViGgFEij7sJOToS7jLHSu8V
6EM0+k8iM8wl98rRRtUrmgqT6lYP/XsiKCl6SLQ7DV8yHIbYnrkfI3bDXx/if6F4Hms/mdMv/m5j
WCqNIkGk+uwIkFQ0cSXCjLHQTC5JZjrRJwgujxmrzcucCvFYnWG+jtDFL3YTUn+XD4lWV0Bscmfy
Lw/BBRbQ8djw1WxT1KRn8wCwFNACxfsVxAT60Fp1T5FDgUjjsbwXAllY6nMCK1P+Tq++dTvh6Qi1
bE10Am6NsoxzZXNMPEiCI5gqIfq5bAI78a+fXhcbm2sr41vXWykXinMzDUAuG4dIAW/Fd8XlF0PU
Y/QTV10n0tHrfOyBSOqC4TpP3Z94wapcWbHTZ75rV2p8HNcqUEhj4fPRNtTQK+pgBdUl80ofuZDi
khghzgp2DY8I8Pbr6JJK+I8kHWtp5xYfecuhenW2jqA+Pn25D+5RsGL2FMfZZT3FbY9GGAuPWyk+
Zi/kRj+tn994D5OZ26w2iM9upwOuPuYyuDxc9wQjI5bkkK0cq0rhMHVmu6pV5rtZ/L8WOanmQ6hB
es/iXpnjdf724ewnvOWXM7pM+T0Ak4P8TAQ5LNUNr2XGiH0JdYFi99ymphTQ1l6DZ7nnnJcjPSa3
J96v8qaqx9uUkV3O6EM7RGivAXieLQ4A9J4N5J1F9B7wEWLVnMF+SZcO8qL5iNXkw5qT+U5iQ9Lh
4xc2r6ONFEEl+bUWiBfRAXcsZttKSFZqCcTAoKEnqvU8JYb9ZSnSEeN+SlCR+iPawXX/McHjMJ+M
D6m6H7TwRrV48KZ2L94GDp078RZBUZbSezm4sZGDMxpjrVwXFV7EZdiTT0dVUDTjoynrkeP2u7do
QQKPVv/43foWP4OuibQU2qZJ7DtTKgr7o+ipbMYMHNHdQt+vs+68rp/atQPAerxjC6f4bRzSKnGp
Jsy6Ocoe6siwBh4Zwxy1UrJrANjVKSyB0HGI1L3C/HC3Ecj9iQDV78pdvrZYCWB8qhR12xYXKUdt
o2aW2aKJLLn7hvH9swa89dCCjF0zOOU9XSmRNKf5hdYiMMNgSDxKikVcyh74ce0uPmP8I84q6VFI
xBoIqHBBg1WeHTOTBN8ilgkw+DgPq53f9oJw40oF8KB3KwVFdjD7rS0Tk/TKYwwGgUh2JxRBwpub
GrMIf7RBXRS0ZaLG7WIqdqNTlN8fklVKk0C04um5y1GU28dTRLLi/316IkJjb1/Y9/BfM6c7TYp7
9kcTA08tmVozRaSMlcWhybxRGx0byVCQ9Hy9nSkJyZ1aVeD4ugARHKXuz6uU5VXGjeqZQhw7BtJW
ufh7cTeIWuzzaxPePeFrOlVXpoposL3k17hjLnC+khLr9BJaT9kjQ8/5ehGPXj33LAdpfQ04++xS
JUz0nLPdhjVdQBmDEFWWV4+fFCoB+RhXZJKsOG68BlTZUPu7mOY8Pcq9WyR0pjj/CrZlKHqCN7SV
piod1LGkIDOBVurrsbFfjXGaOpzdCrH+y2Vdx/3Y6q9cKfCj06riIPPTdsuzpl1K34CtSRQGOoZF
G5viei4HGCOFC7PP9ydEXBIOf5hSkGW6kN7TtEvVquO88Oz03t1EfUcUaSKLHgkFF3W45BXPS2sM
VQcLZrbI84EAKjYOG2GaVQHlBOmBiZNOKXSMVkO963brX5/5jbvVycgUnuhl6QNWMvsq9nXfwmvK
qqdNGbXIu0qdbYFIJ7TXvW7d11pgKxP19Fa9xq/ab/gX1Rgff2bNNHM2yYOng3/cKa1ozkF5GaJX
R5sL19Oycjpqf9bWE/YUi/ogXQL6ggu2fnsVoNvTvvmIcWxVRrrBrfLc7GPpx6tiSJODHxPbLEXw
/5Q5r8q/pWjAK6zfX1OrUKKG57uK1n2VZ0mcia/JLBLdsSLjOCbyP2SaLE7UkwZldyEwri6Lw2CW
4jpWBrmsIrmXsOjbjavRvQ91guEATPSDj41u18zIOlqfkmZMpjQJZ36S6LZC4LayyFBnIwyrHumY
/Pk1PxZs8JEX2wPq7IjetIT68UxJsEGwhhpt07hHrA5vk8rFk41duEk+2YkbaIGq9Z5L83iyBu1y
vE27amelQrGsV+1zAUh3vnhNcPptAet09DM3WZkyxCrcyLdThnw+kehXdJDTWUB8tHTpPHlk7OPY
s7TUpHw1UBvj+3Jd+lztr1YYR8A/l1/zoht8dlhdzXwinSlzEcURPvQroH1kMJHg7e7jDJN8Ahf2
BAeKYG/iYa7ABDvs4+x6kEgsoEE3Na8ZLnIQib3lY5ZVL2k4eIXPn0k9zIXQFm2cfFUTWVDlfkZw
BPSIr+DpdMy5xDP6qOoj8cnEX77JbiVyIdjfv73NtMHSLpv8vIqBc2+3Z7UctaI6pR6yGQnWrAdi
z7WJiTexsqJXjNlP+8qzonK6mZCsYQvnt0MTNeJCJePSppsvPTCyRu6PvKD2JlHCoQfpdhZwwefl
SQ7NqpWZXwTlyGNGESNJcYF2hJ8demYhIyerBl5XpsWIAKPb5+kaWVN84V4OlRb1GXiJxImVeit0
0VaWmunlD/EBUb60b9S4xahxJD5MQ1Uqm3eKy10N2eUXsIiY9PShE7P17RM3TESGrDTkagsUDO9i
MQhI+X7XsQeBgZ6lNu7tS/9AIJVYLflyETHvc9UvuXruzLFcSR9x3njV4nsrSTmCELqrXM2Q5SGZ
/eCp3s5nYdUcszSvXcA4oFW0wyDqtKgV7+mLuvPF/gohXu9q7R/NPZkBqigpXCdiwIwvr361hKOo
nGJW2iTxe1kzy2Fz5ULevd2YCIWa6qUoO7uHfR4LNdVJvcm/9v+8c2ijG8TN1NT4PSaSYLZTwg5C
p/tZycpCOqpk/5tjZiTgnp0Rk1xs2Vcjo44wLKoNDUvKraY2/luyQ4hH2LizmwmY/IBrz2PvjXOj
0Oq133DFz6t1E6e/IQ7epGJ6CQiJSROjOiHm0XN09z+2I5ub/DcfZ+8B1X9nrevDOjKq9/v8W1P1
jRE/OKOujtqR8Mr5n85F8Qb6C11uhDq/JZitDYHEqG8iS159fH8TCsmRCZtj323MrTpeTPJ0jzIa
R49IbFgV+GgY4epe+hTfUi9mKXMQAGaxulre4M/vxs8j2nVL61UP9sdMeITVLIRyMFKSwEatcC6F
8XPuRzYvGOl5Pt1JrKznhvgkc9wnVIsrHC74CNk3FnTA/4X2nMczPFT41NbVkvRMVfKV6ojqGIcP
jy10HD8m4/TFyQzZkbctJYYf2UrzPCt+ePvBAFSU5Rh9vc9qXIhdWE4Qfmpbm22wJTJrlr6h5ixe
9qezcnrC15ILJW4sW+0WP9sJfqUm6aAYaP3AuVnzbPw0AXwEm0R+OK93lzd6223XmxnkmKAv5QDr
YeSQM9ibp6vgq6bSwRhcSeCWc2Zszw0QjXa0bMlJs6tFOfTMGuhYuoKjMUReaLFt4SnE4ABKaP9X
643EYLFmpmUxGO2QPGGS7DL9/Nc3tzezkZ/wU6Za0smgKFq9QuuBQjNkR+FO+/Rkd9qNsWqCwXhA
m9kpilVucFVISFyRGZBDuArz18MKZXkwJjUHwfQoHQC09TDBnDjURZavBcwPLXjFYfg8mnVKeU3h
e/T0WOijZwBJbMG2ZoPytMpSrn4VYtkx2t230J41xteuJ9oBzANZUEMr8RZawypgFDPXehDeNJE3
cIYAtCmha5QjKm0I+CzZWoLu8887omuf4jtutZKhkdKM9kCfnPIeOAm3ssOK2MkckXSa9yebfsX2
1UzUy/6t8QOZnHUBpzGaeEI+txdijR4howQWgqoqpBEeBTW3eljtu4uKAzAqslsol9u8y6ahG1iD
9uQRkwZAAd4Pd6i/2NOALZcS3qLNBTO/0Uz+nmZkwzwFxLYn9mq+ql0sdIuOyxf4iD99Ni3hwAoI
sqYKPQVVW9yv9sjKoBixw0bmiRBy/Wo1P5My1CCqlsTCP+KEPkkOJ4aV8JlvIZsf7l/Ag4f0J/yS
OD2axfNYR5xq+SH0uWpvCVCCssK8q5xNK4AQnrDes8a4RS7Bfs8i9Cheo/A3Ad8Cg1veEPB7ZQr+
CbgBMkbR8bTb1ESa1KlA/0Mwqcr05RYW6d/4O3oEmfz5fk2nYhCpGpYdG28DKX6cuitSFNhh7XHg
CSVX3Of5gI9kmRa8Qong/KfZNtOXahEs91ewO70ll8b1yfHpJ3Vaj8T4dFY7jbJZd1zEvMXRsh2H
ZGfXE/pON2RtOrkCxbDavSRBGs7348pa4Nzb2gSlywdw5LkxtTtmNAlj7hSVzYwPE8f0vVXnsAB9
MLBcaMvJbdEp/WdiOTirYlSWRQmRIthUPFUiYk3KsQELnCORhrZuGFnKO12uaW1axSl8TkzvqiYp
SI56/KkuGEhml16hRq2LnnakH1iyd7/jMBaAbaZXZHSkEcg32uuZDdrFkK4GGIXlQZ+McvXUCkXr
OPeMeFJAofSIl0F7siUKCEMavcGhPLjx8EDSEwHW/dS2TNPAKQkJAbR9VqhSjq2q3p6Wdso9fIQi
xiQ7JlR1uXOE4mUDcVvjK2RBVdG/+/A0r0/bN8CCSz0Jd3uDuq0pMpbIaFPdZ9BrciDVzUuHR7dI
h2U8AwAGJYccQsPnkCDnpmhf+WD6w9wcNXnAvsKinPl/mPtmIagGn6JIYyPFLWq5zOQIMPXfdXsj
sxHR+qpchc/q0u96YAAs2rzH28JEV2oFNIjFrDUTEG0hC6wlku3WhLq4c30HQPWLTNeE4vQZyYHT
ZQUrso49It+2V/INMS8Utm4TiZgYt0MbddEvQFnRSpIgpWySi5ElzIsxwpZHIa9eICFx/EJszfg5
obxKKKg048RyE5CWtpuI655hjAgXguFq/6n3h+s/EYrtGEZCtZcm09ngGDlNiJECCP//hsMXWPK/
ESdzAtcuJqheklQtF1EW83BH0QXjCZyXyeJagdf76zIIApkLEhn1aEvyVi4N6f2XpEUCr3HqZwx1
+224oyU3J9prpCQ4RUm0jlP3fFUFuExkyElCGFa3G2CFLceJWGOKziO56ngZzVEBRsXwdL4tacTO
Phn2JMZfr8Ot/GeIIq7jnpFcneyYPMgg3wINQXm+f9XbYCoP9mgS0ggHIMQe5RbmD8r2L85BkJ1T
Qz0/xjpCCWUcW5CrimFPWjMusQeiTIhgXwCR9CXg+ezxBRxqcYGYed22I3EOMnzamPNsxli5ahvN
all9sPblh9+bEUE4tVUt/8vFiY2NkZzsyOaEaBS9Qy8q6FI14rVU5nvVhpZAMFArNwOOt37AETGH
kLEh6Usm/lHZPhB4h/f7ELHIOMNQELaPhi33FIWEB/e1R85Tb1xSlZDbgEJdkBrhg4R7pZgerW2b
j9I8YdgWIlZFJSyIQnsOdk/qsaCLbpnqSgXEnLlc2hvH6wZ4NuI9lWQYK8JhPr+UgUKaVhrqjTVt
mNtFab/c57XZsK/OmDXOcm84LLnx4Feangw0GmeiXTyPTUJEZCH4OqedL2ly/Jpa1429DNczf8Q1
w9hyMRMzQD9XcU9gfIthYPM+krlV/23jnS4u0sqhj/7CE2IKORLihXfpGYnWN7u0w2MffqVcEGRb
YkbZwYkKlDHIO9+1ZmKXHYioLPCA3oRmG1Locy7wEysIadA3LPTDo+JsL0aptyg+rSToGXBGZJJs
zDkvGLJcUK2gL3hUVW+vf9eNhJwb6aYFD6QLbdbWpVt4E3aGKuxQDIg6+h2OnhRN+JnkzdiHlMj+
SYxY+2Wme9WPDqvrwLbW4AYLAX4fHK8vNwFRtIcb+31j1M6uUg/IN5kYZYddTV5vRo8lKGOg4qFZ
pRAAy2oMllMqOBZ/WkS1AzA2Kzfkb084bTy9bwUFehfr37csV50zThdvJJXWrmYxE9WUa0uoTAQb
Jk/Jrn/HUDa4v5Q7g5E70pkIhoAAFOkpew7/SahluR4DU15uWeKbNjFBx+Hg4Vq0v24VbZddaXbp
w4wJPyNmLECO908SORtvUO6jLT+6xPKdqs8VbqJaSoVzIWM42rZMAWelp2s3gGOFY+1RAgj/YUJK
LAT4p7iCjiilkyeRPBKLlIJj7EMzyOUa9KWJELiFops1SOKYl9vLFGvAgfZxHQdHjFE6FGFDOxRR
/6+4JCh095uRLPpuZyh5r+09QIzsfHcBUCzOZb7SqatOvmyKuIJFOywQB/YkFu8f/1rrzf2C8RlI
siLLkxmyVYKliDnhyhpAP2I0y73bX9hiqV4kKCVapiKFbtaepLJ7gTJolWiXfw2Z9wWIju5k+qHm
OLmWvDeB/22MwvvqkpSj/aBZu7ynxCB6Mj9cv1JkPKdV32vi60hbDOo/18J7RcYEaaMEBPedWgYC
9ukKac8sXKrr7fx88MUN634nCXnyYKjZkkXOCsHgx8S2pNJXc7p3ZZvI1G4doz+NFfge3zXkuHMy
Bjdw60YQrI5mL7eWuSt5CGZaRLQ6SHtsLGrPAgiubylyo6F9iFldyvG0rITLQJiTy4HZYAM7X4nL
MCGuFKB8yh/Z6u2e+GDHHf2SJTl6slH6MHF5dTUNgUozo0yFFYAhmStY1roORUyPxyzf35IGpZ1d
ukXTe3Gt3A4VHBUvjgsOotnFN89Sbea45RdGJg82xXILXBN4o3Y3/nDcsXUBS/1Cv2f2aSx2cGmF
IDchTZJQZd6jbHRSARFlkXp8Ol++kQl8co2U6VcX98Y33qNYbC2TB8I+ce/b3wiSyqL8LEC0OSyY
XtegcKeF2Y1Unf6DuNDUgCvVbEK2nXd0ZlxxR29tIdftGA3NT7s8giuk06DFAH/iV4J5Q6YuQ4D2
669CrBljhopRgEkjaGCjWLIV7R/Am995lIaU5fmgXbHDaw/iHTsG9AF++xereD2XLebPsb+40cEI
XdJ7KrVFmf/e1XWI780daaX0GNcQGHGrAlJSRiCQ3ryW/hpDKO0zoxWF3q1D0/3P+R4yktbT9SA0
3TnENV4eT6vE2f/+ETEeCDB/3PBcs/XSVsFEpVih9xU5VY71eLXey1gnPqv1uj340CNkCE9y1FfD
aOPCx/ps+eKSh20AZi+21P53koET452rtcvoSpak33Gmha1OKtSnjG1WXuvi5jARJsdYqE2g1q5/
LP6iOBsvIYpMew3PxHcYr6K4mSLUP0ep9sAr9rzyGl5lxjwMk5+KYphTm+PQE5HhpfHOTRTTf5zb
pso7KJkiMdXwQZM+A/PNzYluKYZ6mU1JYDRKC++do40L3EYrQr0T0YrkxdHs9He3CdcKFtCGdY9/
qpzDYIU7PTH0Dmd0bGamsZGpLuWS0X50uVhcaRhHSYuBUDItzVNiq7A5uprSi6yErbhUOhnA73ti
X7+JmR9QelbW+eVAkLi2g1ycsT6BaY4Si4403s8Ew/Deu9zbB0z2KhLx6mzD2zWiuIJm1tnZGSOB
OUxZsEU4MMNu7z6IZ9F5OmL1eyvMBLHsmiXLTarFW1VR/5kYBXgSYqlCxhEpJCqmFyblu06OzkM7
3xiAnnYodS9sukLhdFsyd5jUXo3cOXp27jv+WJf7QOW3uaQigqYTjq3FKZZnyiuGLfkKq7M8fZ+E
+cWUoT21rppupWcZZfghuhxTdnfKy71gbD103iaFQa7K6bqSBe/pELy9NgQeX12g53xoh4C32zAk
I/kyDueQYTSpZ0DGvn9yoDzzV72OQc+VVHkO1sqdnW/9SZjExY5toJcN5j7qzUEcfnyJD5h0ttvz
YatuR/93oZYgLx2aOMLJxWzXRViK8BvwZsRuFj0FQupwUn0x3N6pzx6HyZ95s15PWycCTkzUVnuc
0jBqVz2EUiTzWynkzoDvvuPc323yYnUvmmwJvclGa5ziYWIIxfB2eckPgNhZY1muHgJGGhmwydo0
GWOIGB9mG4zS6/zO7R2yib2H+oMIKbGpMXOKo6ZL7cCSxVzVNpmiEyDShCDIaAuedrrplk8cRsfI
QOJRW6m2fZADvODnVjNl2pH4myYiOuNn4gbOEAk+Xx0943cPs0LF/Oin4hHSnfqfeve+1uGZdjiK
nHf8mF6ZibuA6lbb/UgQjbZNmJQrVJ7+FHjipmG6ExKJB3D1oF0QouQkeyTv8hmY3CWL8K4cgNhW
w3L3EoARJddfxqJo3KKD0+eo3y7hx/jtgBw0NwaEUmIkJEVF0M/q2Rev+IaJbnbLQKvukgxAKTxF
iIk4NnMm9XvDfr1dJ+H0eAcZHJEffNaPAQvoqd/FZYrzH6LMbjWsE2YJ4AIfSzCDMG0vC1P4tAew
NVLy26KV7epgSMSfx0f9v5tCJ+jOBoSt5ZoSUR+3ieN1icgiqhfa2nsC5Dl7UUxMPj7I/4c3KSsY
Hxwq0xSkTx3SpgU9LCOezGq0I91ZHwU5a9PMtqhnZQHx28K8AxmbANSjBJiIYvvdTL3EdgrdPiON
Q5JaouyYwLu8r55MuQYh2uWWBrrA2o+S3f+wC8NxXZJDRrPh1NKs5tK9mbIBvH3QmZc2Z9up2VJb
hB6WfO0P9hZWoiDs1C+nSGuB+6vDKZMrE36nqT6uc7du6j2hg0URyApNLGXbn3lkGAK1Hqbkd29p
+hdxzqeNgzkH9/L3wIap86vwX8CIbpAkrPm5XgTs6TNsCiwWKMBy2F6Hio4L75bPol2mGsHen3mP
kyM/MYPKMJ6J58EFmheZ7pzWffTlReGZhr6eYHyf2yjO2N7PN+fU+FNXvO0tR3sLz3LkPlml73ZY
ws5x0rs31VwuZ6nZ81OF9q7ETwu2lxkagG1Av0/7YlH24U+QH1ivlv8uK00Vriejdi6R1PinPYgH
28NQAwY1fXXyPmBvQr7B8FzvUPrM4TdGsHbvL2xtTx2TL9+2PGJIFJV52D/TEHcN+x7kHRTp2+su
3mqo0I/bE3Ko1qkfXysQV2UpcFletvLn5kO/QgZCVUnvWG8Zwfm7uMxsEFEq+KDZopKuVanOsmXA
YnYby9Qe9oy77NT4R5fP/oy+9sqyoy5nrRvlV2Jn1/UwnAKd7fKynRv0OPtXB1Zc0zM6zM89TMTJ
emVGcyxH7zUtRUJdt+5TW1xDmExTTFx6KkBLg8sFgqn42htrj/V6VpY1++rRl3QjM2OSSCq/se3X
60WmpWOCiyWZXvXGJGAYbOmoWPxBbf6yQhDNXVqYl78QF+DnOyIgbgKTwYNWEwGTNfw7Xo0WM0Ul
dizocsREj5TtiPSR+X7NdJ8UID7WGltYBvPy/moXLAYi//M7kwJi5Du6rdjmO1wVfawisQd/TEeL
FBo5oZ/KAD0jTU9j/koRv82N3eGQNMCRZ1XIPO1cATh/oR5H1R+AJYNJs1E9koftIwvTN0uJ941L
5i6SnwrEodbwrfJTTQeg1tMmPbfh6aSRFsUJEyt5gZGrmpPiXT2byM7zzYiQ9TZEXAKrYG06yjrN
BfSWUg4QmD/ucj13OlG7nnmR885TEZMCGi4MQfm+tV0C5peEJ2qBzSS01PI5MyOjHp3s60kONOoa
LagrgRqv5hn8cI4oIy8a01yn/LJF7QDWSzs4mkU0B2PytX6BJQsQMzvOoHY0tWzMMOxP6Roz1VnP
s776/njL0t28x/BVSW0ML59zvvY0sLxoCI9PGh2z24tYYcBcIEu2QZKb/uDWQYXRzSufcoN+mwe5
tZCdnzysbCjQAbzjWJyQBk3VgquL26Glz6ysDC5Fh64zX1hOQErO/FpPYGkTUB03IwNL3jtokHce
ZPuKDWevI+PkzQ5M7q+QQQ/FPJR03GGMfOU7wCIUkUDokjZIepAl4YyyryXhqUH2Lm08WKYjNc8X
ttIyMIe8NgByHF4w2+IlJPbEhic55UP35naJ7WNAa7hhIp69GqfKr/SJIIJgB8e8Jy1jbQd/13i4
NI8Q3mAFxmsJGECWA48JCvqqg2xx6bkw3o1R17f40GmaaGVYc+4yQIWk8lXlVxLRdp8wnw2BvhZ9
n9EkT258/YYUmMyOBys9spKWXgTEwU9D2FOu3j+kiVFMtrwLYg7uLT56hdf+udONA7ooRhjhtqQI
VWlA3jWSzKssi/QTnJRk7aNuMGQPEOWDrpgOZwP6PXhV70QeRD2PsLtpk0suJ0ySImXDpRNEfFtJ
lAVCSgUIO6U0H2q+ztna3aEGUJT4TAjwbfSEgzDdMgxzUaLfoHFzYg4jMzIcVVMFBzWNA1wAWhQJ
SY7/aEMe3TbV+alsgEewtcVhBH5MiUrx3YUq2B3kS857AT0kBEkJDi0c7Z164os9eA+ucUPx5c3r
mKUpgJ2d7IiHOtf8sfmkoQRCp5c1CXvJeFgpmJZUm872pQkzidqO0ixgJzoCuB6XflupnxCtXmsf
FWj0jIOAI8GsfHb2bgDgNxSfhVBeSdzapRVMXVm6oWjhC25a3DxLnwR0YLjQUNJ+8BRh9cVsH/cW
PMSNXJwQ6HY9kpdCseDAQd8pEzaXh3vs1xeZYdlQpD2s7pMX7U2xLqdbJEPV4PcAroQkDKyz/pEl
0DRYMnJOFi9s0HDcrH526s9x7ah2abfeXI/EOHINR9Os0eGhlQJ66TAtrrnqoxSQG22vrCpF5dKM
coLoavzkp6zHLYipwuE9BsdaRuADJrHW/nUEl7l9jg6guuhCP0ud49zGH96VbDWd5+Xs/2lFHVfB
p7dkotyYBQHwWoXe4CkzL5n9s4Wl/L6nN1yYPpTsRFn54E1fvco48T6iNcn6hZP8qPss93tCovk5
SOnmEH0YV9376H2vgd0LB97M5AZ5RNhXIzNI6s3jRI63HIi6xNJfmPSJ1BJOGSAuHlaZh+FS10WH
JG6EszH2jm0+Kp5R1gQbLepwTX/QrdRORsn587slHnkK7uxrf2oDd8084aXcO2oWQ86iqZjO70fo
nBjioanZQBRZluispVlh/Xo8yY1FrLquZXH806E5eQ5fWAXV/OtuhvX1J/QeR2vyWtoZRbmd7DdM
NqLHYFIRKmhucT8tu7iRcHwcda61XUXuaXJwIZsDeKQQBhG6IOif9chSVReiZ8uE0hJN2BSD3yVx
Uqn1ExucRea4t8Xox/pzytk1NGkT3Serx250zJkzq2OCMEP17IEGjEEpOBfdbTatJJWrf83FE7Kn
d1ECpZw1pBpshDlj4ZFL1XuMZXYaNQdsTYja0vKecsUjb9vwSG2tzdwJ8MmJTHgRl9FKNnUzUeIK
sTFgDJrfylGHpTy962UZN8JEsAPugOnr8IyA+WO+PewMCi2MKoDfePirr7N2N7eLLRd1gu9Z4Xez
C/uoTWPrfPCvQAN6ke8MipMNLqfb+rtE1evbby/oqwtLM22lKMKYl/w900nj8pQIjr8garsAzCDU
YYcImQBu5FH08DMhrxe44CqyeFSoFdxf4k9ChFTtup5I/AWldLHmwfd3jm6JeGREX6H5bxYZTTmT
B/toRo1QQ1qJFQipfoMmEAC7AkqYyPoihZGIDHzrqI+5d+YZCz7SFB9O37gnNvZOKMzT9YnO1kWj
4fgdKsjJp1dxTT8hibtzkO8GPHkvY6/zvgcy8s53PiWYPTAcH2399mj4BbvnMcWcXmA1D8rxwsO8
0jX9jGk53H4+C+FlCStxoj/pG0f6a8tQf48RhccuBIoYi7T2oabxEdRKYEEneinfBSOzwbgOUc08
13S9C7IYNpMGOUUi3rJyfyvFS0Yxc7amk/W3F/a1OkzO/n1F/7gwCYwh3yyEscLwjq6hiVmwcCit
zuN3Ipiaf1vP10mZgf4umzLu20jDsN2GavRBtoDVzyMPX0LRno7xNftyMOiCdO6eLFhdB+kAk41B
qq6bIKWVgwIPh0wIp1t9xy0UZmGXePGXt3IeruynuetCX6OqwK40wDv18/1ky13vhEY7aIgOfbr9
sjmr/gJciAshZzNb0OFfBk0acA2sdDxo8lMYtxui6jzItR/cosnbILJGbrtLn0g+dWwRQl7xjmB4
tUp6QCDHckVzsp1wGslgh4b1fAMWIq3B7VEY980v9Ggi5tWYhRuY1vmB7LmwHId9TcQm13zd/+/+
vjJTD6BHlgiqmUvUxPZJPCgdvKBX0awA7ZpWZou2uAC1ovDJxYRcWqPiXxFwTj4KoM0YwAhE4kDb
rUuOupEuIg2QzNM7ZPjYw5nbnpmZSnRdOavH2L9rh97XPyABfISuWuThdLL+QMGhrMmmNFizROvn
XIfoNeo/Sp4mOAYG3kU8n57ugkR+gKfyM88lhw9wlmc4YXGDBdBrv+xciqYtJzyuhlfj1D8Iet0a
skHIaTnvV8sXHvSIHY2glIncKHFRkI7+3OlRgXh3fUDzzUSlyYTzp2SgVFB/P/pCsEEaobYu8rwH
8BUlZF7ckFeudqAze/TL00od9slrDAf3sanCVZGE0kx4H6hckgTiq9RTULRv+sNEMuf8odazG+Jp
Ef8ipVA3Fw9wJvGKp9FrDijO6N5WVv/AJgnhlv1rDqKElzqhRXi/0StHD5o/8wAF09sd4b9Njhyh
bUzfdAFKsqARVlphzOJPIdTjNQV+ZTl0F6AN8xp6WDYRJRE8lwRQwZ97niUdlP7G3g1b1CL+MC/Z
W2NDvdT/LZOL/az6AqQjOheN3CHWzOt9L0eZD/1B89SpFHNUZOYEmfed/Ki5Cv+5WEZIyGsevxqV
lmmQsYHBM9PS0q8Hptufrcgr1pU/Ua72Pgxz1A8LdlvLREJ4ygcBEmBQidDokxxaMMhesv7Ngm+1
1TyBZl+00Fvb7YHf/V4sygXwexE/LqEunyx3u6f7gqJWy4Jf5sOhpuRfotIbb/QqVtt16gsX9B67
zw/Ieh/O+7/PfPGZoijp+A6TUxpLLvbqKZGggmYzoLglTrwNH8gHONjsKX/fCbN/+I2gloUPhiX9
Fs0613GOBN0KEh1l9QhTBVLvda4iPTynwvCrNDAFV+q+XUL8HxdA2L6O45LAmaiJvfm3Oxccn1W1
p+TELG1ejP4tZNvQXdifxHr27cufqfjOw3w7QBd1CY32+bIw9hgmiyzWxOsrQYDDLyHrfYRv5DAy
h+YaPlXBpR7g2Stduy/mzr6Qt+RlNJ6PqEQpVCtMwsO9tTDUn8GOYQonJc6KJc1fsde583R65b5h
uAcuR6IS2djvxsuHYp4xMMt1tRN5ligBmOcddIx7MsISaf2LSav+lis7aZ4YNLnGkYbcFP9usOG8
TmTOeuiGta9poNPIuodQanlyoWJzzHE1KWDpcI521kvZb8Ea7uK3lo/mTjR3rPE3Y2A1MXsvl2Zs
IOI6HnpkbGNLe57P7Ii6LlzZQunH0h/r7TNlA+UgOSELxi0XEFxsjjVT1Ht9Wtuz2DrIWd7wlIFb
ljxlvrsBxljOtgX3eMk+WtHmJgZkIJq3cBJMqhi8y6iZF4pmeQ0JAOkBxtpac5FeYMoEPvEN18yC
0yD9dwCBweQlbkjWUXjj97gLwLZHM0/yF9qvoAVpFW7XDhQ8yx49eHlC92K3+VFrzXdeCyE81HZP
WLnJC7I8wzp6jcMqkC2V5CxsQyoNG7dGxF10aqvJxEoZvCqqm7gupMZEcrzPT6ae2kEkYvR5+GUC
YEsBXx7WpEARkJkss8UhWdYz2KETfaUWauvVkovzMEEJvJq5deet/zkyC7vaZdhRKmpoOMCCQeJQ
JEbk7akhXc6Bhae87yOWbnehcOhbMCHBMJPBXWX9pT1fHYbAJi910wotRty08tuPWnBOuhqCIZex
pWAkzc5gZUiYexycHEtp3Q6n5FAQniQRYcauTn9Rh4EvcqR64yBXLwFY/4PAmWXq0g++7ZDcEK2A
xV1fDBhY+Q9xjo5zJT76ljpdBZaqUlVWxph6rxXblKeFtqxdpngv4oQtsRu+xHCPdaGab8SdrFpA
Knb527ls4OHKlmjFObVSBhBjCYpZ/a4MMe3FPiKvOef0sxaRXhJJ25ziGuH9IB3iwVoJVz9Ml2iz
fo/fu+k0bGl7GZad2ifJrJsd0BA8QGbBfxCsqNyC1FK8NKQ423WXDT4blsnwU9ciTu6M4NYDPO8e
RZUz+XEUXEENv6DTz20t5lGifz7YPrzV2JtV31o9WIhznxGNldbwPU3/FM6xIZ8iMBtVAMDHSauM
E1tE8FQXOs0jBYIpGBqtWalz1Jq3hEubdAQGmglkmGgoNUODf9rE0wj0F6BuFhiYK5WsnarhOk6s
m0xlX6MOt/3R9o5g0fKKZ49QpSpkbVj9ToChXClyptQ94fHc51eze3y7Mr7mBotagQFWja69R7GF
6/Aof3gcegOSMm9NusBqCSoeXdgpAnZL4XuJIicfI16meoChxIT+zjdBUqLhpVxvYgQ605aOnsez
GJizHOeiO5LoViXtRMsA18XgHEnxZrioTixJNkLX8PWP8Ur7296OrUzkyPE6X9cuhbjQEqTZdNQQ
Kr8wcPGtHgkh+xCfaAMvK89gfZWNGt26zd0CGJWoQbvdpVqSy8Lq3IdwIyyVWkj694/dPxeuVEX/
eRkEfUNDvgFPQtA0ebquyOorQSoMnc9i52pbp6WWqG7wEBCB4csxwbM3nGoYOkfqHO/kieqFz+VD
duKFM3QOzqrf5Vyzsv0sK99fpAulB7K3NgjdzyAdOwHx7l8ZJGcCTf3dLrwAKo7k5XxgqJ2zf3s6
vkoV6uHJZbtnXAC8KHThw0q3XUTAxvKN6gJJp+0wRRU0EU/5DURexwgsEvOxI9bheEhjvfNp7yqq
mT8Y9kPJs5zYyOiQCBovlRzocTBwlVHCP3pvV0KvF8s1RnaCFBUxnVZDQfEawk0bgD+E9c15Ovja
xjdk+zIe5RKnV8iR1S2D1qPUqtDGTxTltgFnbj3QX5hABnb5hJk94eoyV3y9wE4FZsRXhfyHgNui
VJ/JsIcTo/zPrdPqwbOTS9ODEW8ALrMednYBqn12HmtrQCXcZuavATmzB6Qw6ZRWcevunLfOKdBg
U8Zzlh4dbTZHlLqIZn6JEvC541mLrKwK7SHuaSF++nHNutc781MHRJIp6kX0IUtkp8yIcX+jtKna
bhSQvdofYMwAYbJRWljtGqt5br7uizqm2btVm+M3rhpwgxh4DuU+H/chpgp2Xo9Tdk8LYs2ArFUw
jR08k+vB1fwaST0k0r5+8nZfgxbbrdaudyqDatU2L5rgaUo2xQ0D4LsS9z12lKGZJWxnwB3CtyTl
uEPoEwrkUTIUSQNktQ4jBrH1T09SDRQIr2xXeZ2AgpqvWtzs1LWHkoJnQ6alIfRC+jFuSofqyl3J
Qc6GHWOf2lfxq8+x94Ki8194W4QUG9krcmulcA2R+OXmAfqov/n6zxyXYaSmQLu6acPOhYQaJ9i2
aGhPVOl3zybNFYUmS9ETbeg6qyzQlS79ikWbGXbV8jBTkq2yGf4y0s0jkN6LQRIP7RJzy2T8jE8v
eYJNgztFUvFL7QcxDOZLZgyw8Pg/H/VVORil2tvvJ+LheIZjnfaM6sqNPsSBl/exjFpD9yxbJqPx
rVsHERPSmcq2QPD09/YENA+XFf0FLq54X/JWC2uIV1RpUkKBjwBK0VnNOMZelkz7AktKRWO1CW3H
Vcduv8rVwvgmh8liMZSnG3S5CcAoxyv2MDZvlDuH8BSqHOIET5CMs8AAGMe2vzPCxfi8S0fnJEI+
1DUfXwel9ez323IUzbVj2UrE8JI0ItUJRohCBaAvNS3zozFKiMSf3BCgBi0zEZt4rckLVElGTSFy
LhAS6t1Omm26GkmF/1x4pKqaaiO2lxXcrhsWQscajId2LJfFFkShGQ6ioPg6/xXpyW+2W0WK0ncB
qwKUvl2z91c8n/+aQkMg0I9hzu0qluzLSPv7aMUb34fmVKXLMHnt3jC08YJ/ju0yWs/9iOFvqtN+
eqBU+7IEQc/vR2JLuz33ME13BHaV6NKJqf0SXZ1r/rHPGYiH0LJ1CruezwLNYyb7GgUf2h1bt0ZH
viYdjlFh5QGnyfr/NkJsB6TzqzWZyOyMEK9R8PbGp4rr78TSal1gbPIflSSWAO3pohBewYs2ld56
jW2gJESrS/mTpImIAJETzo8jUBY2X9QzG53Hjm4ynwYx1RvV/hv2y3/EI6HIg1JuuUOY110V7M/g
NB0i6CIrBvHL/J6sKPNUX1BePwDlirRRhOzJif+eKBk6ufSSR5bzSdTbJWYphyAlNGnbQx+m0CwM
WU7AEkEcZtgVrDQSt6Ee+rHGhvTVjzEatxg+H0iKHb9JA75aQI7bq5WIiIvJabqyAQfi9LDD54Rk
wgKUQqDewrbWdOyAr9JVDWlD5tn84kfeHNJqprsDkk6O12kLPSau5aOh2IUMfoU2Tw8rMDuqEEwY
J4n6l/1WV2+vu5UoNtsJb4/NBwjGshUu0M70CQ7gWfRwc9v45XwcIfvusebG6XZSuYKHvCJA+v+C
y5eN/26s0nMBliAdaSp2yDHBemm/4c4zawsaWtniOCZGonvRU1vYgjlsEOIYymhaQxUHZQFCelzz
g37Wxe0gzZPYVxS5bGME4f26hxtudVhL9TQrQCp1vfvz1Qz4aAUjLRih8/3MjOpL+qqYoBjDevkB
6tpPrJZNVXWe62I/05y6UZ4wB/s2lIVg3pEPb3F3Xs98Tvrk1lMvMQzQYeMuw+6HgECIJFzxCDGr
cOFHiOJpjd+t2r81rlcurra6yG2LLA64B+lShEWihRO3LhZSsSs+1L17v1AYBthdDr+GbhNBD+lF
QfillNvTsLcDke8a7s3YSQKItqDP9Pd2LNHyBjVHmx1Xz+9U/rISPUpKwURw4VLUihj7D8FYCGdj
kaA1piDnwTm+pSP+/h/weI/rOL4vWSfvtaJkNaq1LHVhpOFWWrRCJ2Wfxx0Xqgvgm7bTAdqLlT3C
5bot+N2Y9HG7PeVyErlzo+FkbSQxfHOyri0O5li07ta4Ikh7xtZAP/x7mA5h9U15+iy1MxsZZAal
SqhlvR7FEzGxY9IEqdEqwWAyFfyjBFnOJoJLeUtt58gS/Tmb3S+vsBKnOXJpmcoXZbDKDwOy7Ffw
LfBCKtvMZ7kPrazDxPHmwb/aAbSYSWysOAOFsVPLfAdBbbvEId3occT6W8KXdgiucQ0w0SYdRerc
BsARmpGNivrBya1iYkuMGdp0ZphcSFLxQhUSWMGE22a/Rvr7wKVUVgRA9Tm0c62mJXquDrd1Uzl+
bPalhf0kL5Rk3jz8pIsw0QEegnl9MkIJ3QTCihHgEOrGbiseN1TlxrBjD7oPE++Vu+jgd8A4gK//
wwELbSQeBmrIMc1uzVI/AH7ThdterSb+/bmm36Lu59bRzbqL1phohlu+2/rCtx6qOIrHFgo44Ob7
qk2PeL8JE6lZYj+/FNAnZJ4cqcl5aJqhfM6gxJU4DcIB2R5rRGhhH7WoNRcp/kTEm0BYYFkkzDP8
WIl1bSXjkKJay9MKVLKkXBvqlPy5qIdlt4oWrFBivlRR1SotVrQM9auVUgAYMj9u03ETaDsb9Hbh
JkrxVeF1cuR8cSpqnwWvNp54jReK1tk735PumF05bRCMt2i6TKZYmxMiVV6IxhoVV/t2EqBlQ+aJ
NxXCzZznpZstz7xoa6TtcXrGwU8aOpE+KyRojxoYT10SOGtQ+4XncgGDuM4O5TqpOLkL01uir1/2
nO4PIFTrMNTtO9vj1ytKFywtX/H+da9PnolD2P95IvToqcSpeEj4g85x4oo7Eec2e4Lx39kB7RvW
wG2TWraATGnnr0KLljVlD1PNOkhwt24WgC5BgTw0IQdrcXTzfMqRkgdo7USaqeN906A+LZD1lTFv
nQexczEH28SMuUoBMJHiVg6ruAsqyHnLC/PNLTjrE/h1uDsPr3sFZglDOJ6F+vqM0O3uJn0tUIoE
RBEckzOXdgxQviH/K39PZUoJIXhiwowQDMnU18RAxB/rnejaTnak5ygVT/C45WZ5yLC+wRbOhepX
bRpE/w5AL5dBlSPAnq98fK/3FmdNfy9iTkDiJfdUHxAQFM1mtxyTmbJh9Zj+j0ypOduCtZQdeRaG
QAgK29Yd0+jeU7VNXZ6kT8JczbQM70HIjbM3vH+e9sFWA08L/72FJvtasy+9XZRall9ozrvdGsCs
Gr1azRNJXMsNGHHFhzjKD8CnicAXkLvJ/iE1CbFCiZVNKDFODVUeoTnUGPRihd+VzBW0EOEXNVLe
NT/e/Pup1qv0IbyDFwdX9s/1hRyFaCzhgWrR7J7HEwmpifXVS93We1duz+6sDZ+/hP18XY2xXy9N
p1TJ+LkzVorj9Re9c22oSll5XBmKevu6NNtW2RAdYDeBi7fgEkmgjoOonFB/WrSC+oYVADkV2GOJ
8uiLUId3DIhT+J7+I59mjwXQVVK/zPokXfKvF/ypier+5p2weG55c6HgtHNIMo2B4lgYGQbRykt+
EMZpTKcf7FTduCBzXj8n6WQ4chJsP6kUBZYYLksLw8XbyeZwZwNnIos/FYRcPqRbTuJkBccq3m7Y
cggdEf6MVjyoXEO9wNu/Bgtq/AKaA1xCBNZVjRz6Dlww4tzQ2wrVaYFQzWHR3OSAARPOg1q+Wccz
06R0st/grkL2JCYeLOw8rndLqR2BKHGjzWeGmpK3L2B2A1d52X7SiwXUjouvi7wUNVmTzjbhRdR2
inPoKQsx0XzL1XgfOF2t1GAr0hiTCQK8//pVC4+AAouYxgjOTE+TKhpl1zgTcNOzuX2HGPV8IIKo
8BQpkQrbP+lAT0jGJ5Ylt0eBm0LGr0yvbyMxLLrIbn/6evXubT+fAim8xkS2O6hkvj1rJKPP56DC
pKZaDLKg+vPaPwepTPEAln1VJOqGU8bPypV89+nW4xUuvGW/tojq7ojUQCl1eXw2odMGBpp+X1Oi
dhCM6ir2kfpN5c4lxJ7sSloDeNjlYgGDjOygUzDq3+FAtmVJmkPNPZN6zUozuBXWDc2XOG2oF0ip
YaoqeiXGD3a1/IY7zIDUnUfHAqKZHgN5BIBpakZi+j6q8c4E4syhww9eSKSLkAbFDIt4D85hZ6cV
/MfED+fZ0qM8feCIVOdObt4GVvJFNLjzKSCZxFSh+vpHeoQQr26GPWAI1hXLmv5rwD1sAcskGYfY
B5lyWFstmmt/S3HkMycsSyzZcWixIXZscU9Q0F7wvroETaOHa8isTzER4UhbRYlcuW7SSEBxuOXW
TkHWgKPr09MsoG3e299gp0PzrMZPtALVmfQxxD5cP4bERRzlh2HoUKdnTGnRtyYOlvRxgg4qWliC
nVuc/x2OKg0e2IcJTTh6R5qYku+/aAMnCvN90HUtTEj1p4kSoUu8nN+krBn/NxHfPs9uBzWtyfC0
fW1sIegJ0wCyhGcW7PlxOkTKzZmUJ71z9ANGsBSzN9PZTY8+/N2jfQSqF+KoLc8VG+8ddXYbkOsI
G+3THWxyHEVi4BDeglGL6i7FdJmvlTwtwKLE/q/rIq9iDEmEjILTYVYGxQpi9pgjO3/lxx6fJuhS
SMMGCAHoE7fve8XnG3PLjPq/s55f9ohYJ9mle3xSJ9r1WMEFewfRXOLc4MojY9HEEEcW4JqZWOWR
0pYGkqjycjHY9Epw8hWJ45XRutnoVjjLb8/AAsoEvY9LVYbYolR5wXDF/NPgBZeWugV34Md8Dw8R
W3t+rlB7jprauYQql9vkQV/eGmqYPpOlQ0UMUEEtmP5+IVlNrnv6pa5KMOMERZyt6oKEs8HizbP9
m4oOl8rKcK/sxwpfgtq5jNSYspLvKPDGhQYWdpdQCHmeGm6CSIBzzY01tQfztMu/MxmWyNCd4nVK
teBXm0VN+he1VvuiZfzM4gmAHnBWWdkT/2bzEmtitpDLhj/2HkAuoqPN6mKn9I7eVz6IykF+4J4W
pFtzN00bpldUqqDciv0ofnJZx5zDezs+Zk7JmSlevDMTKuGakX1TS2Q7uta3YahYaG/aB/BVD7BR
xIp4crU8uf7XYzxLCdrGhbK9zWtPpSo4745Zvmod8OKymt7oqI/M2wFPlRJhSDboO/X97yNlseka
jLr9CNEwZEs7YSh/PfIXIK6gYDXeJTgXqYEbcC9GvecUUA9JjFUBvZ54XYdt0/sD4mZ6enkJJAqd
reppAm1mHgkqj+ae2BTTUQKZ0xMx+oZ6mqIfoCXOO7C35ZycN/JFd5JWlcvWQcBUFC8KNIeW8JO9
Ih29addOxn0qvzs0a8cF+dj+SWwOwuLU+tO7Q6wN5bZc8GyqqH9onyQHo49DRmgeZ+KSWReDlh+x
pRICARyRYTYWBG5FqnNT71nzmexROB7cymtoZbge9Eawnn9Ft258E3NLInu1aNS67Y5JpQB7+TXJ
69TtTOAeB6MfkXFjjfQTJGU04rDXikz8TWrkkuYVELAROeExozwpKtZxGcJd/2heSi6uh+KhHEEz
odujCeP2lKfM6fwi92CC3ppXk9puTZ/4AFCGA4p/iehl12tzwweaZKeddSM08n17ZGUCIjS6WdKn
BKq4NF3Y4oesR+rLyR8ZvbhfGMYrcf5xo3zKwhTgaS+HLvbe8GH8/2vPeAKOYpooc30ktaA53RMa
sJGYOiP+W/+R94Hx3zGAlxw17wAQgTnGpBBf4ohQtzfqAn2iLqMBziUlrUWf9tn/M4xizLfUF6ls
yIUmN4Xhp9yOB+SVOmfvjmPV7hdh2jiSKsnaD86flACaPGZxv5zDazLQVwGE+JdQCbItkdKsj+ba
PCAqtftigQMUV/PkC0kHdJ3rCJpYusMO5MP0N4La6HEk2/BAJt6qHSIia6gN4Pr7kLgeVTvL0BdS
bQHrzG5P4Bp1AwxW1+EpJulfeIgw9ab6NDChYKSsHGcgk0+3gRt5Krz9bGZFKWxwW3Qe4VsFzB1M
myC3nF55zzTcQTmwuSb7KuSs07Dtjw3q7Gx17xSE7ziIsZbeRKzxPs4HoIvHVRfceUC+GUYqSqY7
iHjBfhxZC105q56bcxHu++dPdz6wedVV5tUNE+gjkxhpnRVVaG6aenqx9CLb2w0AIOImF94wsmSX
GZYHMOw40IYvMCRxFODZRii6y0w6LwSkLzFM/1vVvSsFHECtDWjLkgN0AS54/fpqAXx79DL+NG23
8KOLMIeKYWLZr4JHe7awmXul9XaZqIGlZ4aW+WADeZM8Kjx5o4GOJl668qTt4litd8ygwBusiLiX
TB20/3XpuAqEIvwX1CVXhAXdgA4077rb4jdjGRumpzchew54rS5wWU2Ztw0s0ewVXKAxXk4I480Q
Pffn+XmH5DOCleVyttnQCFD8UazLmKutiFDWSUHJwmUViASIaoBSIJjm24n4j23Irx1f70c+bvSe
4wxv8pJofGhnXDmzazZtSf9qb3++rw+/jMQhTPVubFECMzDYv7HcIrZy5hxY5HeLGo8Ymf/fe1FT
1ppl5GXCz5Koco/dlE2Q2IxsJt5ZOokOOYo+P/SIgRYvnAVTB54+4zael76aQ+7egtBXaGSWHGyQ
stDkw74cVRQ/tlxglPlqTztgNm0hSeCJLzagbmqM3KlLlyciavtQOGXEsIfjoTFL2NUHsCoOtHyN
mg3v2iBNy1+5HnhfX4bgdHmyCNAOh8UofOXuSvlDSe6LPPXLV4a7bJOahAslk+2cD1qBtNnuVNt+
qm4UHUP9u3iKTxFBy9glyl2smvLIN2r0qrTT1zPsaLx1hrtVHvpNDdnnPxF6pEV7hjWDyztbtm9I
P2qNX6scRcMzd+xUij517PdCbW3lhjVAw4aqo+d3hJqUM8xdCnx2plZayaLrktoRCzJANSoLsxIw
9K9+5bbx7vOSmDwFufWS+LMD9sd9X8BLBpFNL/bO0rqIOdjB2Q0ibeFeoLPg1F4a80cmG0nCzmnt
aeerLmAPbSw+S4GlSVRke+PlexH0UUAE/aKRR/sVgNofaRjXp+v+eiH9jOErOgH2Qo4yJijzt3cE
7czxOoNGcMZaO94nTbUMjmltHDhF1Fa/htY5XjSQn4CV2KAWZmhV62PP0afAhun0jUJnYTeatIsY
n3Db6mAGVqAy34pUW6gghBv7mVrPBr8IJuV9F/vtS+/kz/YkwlvvGYbm0R4nJsRfdgsteSRB23+p
U01iRmkDN7rCGRy1mYJ+HIRe2o3NPM8F4li2wmGW1b7Wz1KfH1j7uo250SOwr89wS47HWE2QgBZK
/mn3+xHyFNvyIuvYZ4IC6aYUa4LDJ3QWCXu4Wr0RFQaQIdVwJ2oKI4PLp2HULmMNBYNEuGgaiZQG
15xCj2EdOf/rQZdxSpek/o/zI7N6wlTgjV+vrAW3Q0sQ53bGeBXLdd693g7fNJUTMxco6/2b+YRl
2qdj4WTVJ+I5ZG2m8efDdG1VLwJHDd4tveAzw+Xqi2mqKPWpe9FbTbCqCHMwA2zfcPl55bNZKpMx
2385thFvWoAtPTTdQGUS6a5bbaDWddvnu+p82OAub+1Ozojksv7D7su9kahlX+55AYwLU8Ypdmmx
tWxdcHUpHzogdRMv1ewtu3Pe7piFGsNZ/i44htOFhN0E20Z/ZwdjWkIspHPtlGZBsewa1smJ68/e
sfp3ndxP0gm/v1QdiwIX1g0SmOJPVCSbx3O8jqXPgbfExpgabcgM+siQ4DeCytWZdiIHMV5BLMx5
9qbQE5Gt2tZIZPvulix72WayyAd/5Q6yYuG4rt8ddFz6MpmY7FJ9LqYdxawX/2UJS+cOgE5XVDrT
HTObjbU9FdbLMN/sFnQ5XdKpojsNQ/sMGRLStnWDWcz9LV2c5o571dQtuURiuiwmeupABr/X9FoR
eBgEOq3i7lkeV0hcG7MvO3hOb0F+O5vr6rEH3NTqV6D0zI5NhNMg0O1OF5N/5fmcwSrbTOTgFdVp
Zso7Bc7YtsG7IRmECJALz5xFdtWRJreNIjJ3CQD4y3J0442rWeYpc/2qYQiHC7dFg8WcASrYJR3q
S6ZqfdbNpyvd1jZC8JRzhZ4OZpV9MwcVAG/+0iclkwc1K+pyXwbBZv+rxSi7lAf2qjLIAcpC/VoT
p8tKbX/bnEM1iV5ys26uTRprTqbosZmqAc6jQzkFQIRzvsRPRMMujxa86TZkUDUEre/YvfterC7C
fBIPqErJYc4qDYlm+twj4WoyJLwPuGW/SkNXhsoIAsbq+kAC5mjM68aALPC6hRbUcLLp8J6ktp8f
mUd2mi9vtMrTlKfZ7NluLjs84UZAznNx+HXkeWWTj9XJoFnokbg/L9b6kMjnZjkm3KaX4hdXiYGB
Lcmag4R6TlOPNgh81dWS3Yohn96IHPHNl+K0WS74SO6rv8USeMa2tO61udrauuFrOsV9EcsBKpor
fNThS00eqhbEnR4ZdJ1s/+TLGEhmJjwyDXtps116v6TMeGBXSQ9sqb5OdOvZF8jb51bICcEE9dLB
DGqwW5tDI7Y7r6IPCTVmYbtjDFeCSC4+mH90Hv2trMQ5D9HUk+S+ZNtFpQga8w0lwHbGPkUCLJPI
Zx1WmTbjn65AP4RxXV7+f9uSWZnZ7UrUu/3goM1225db8XD+mq7L7TqsAuuKk5gt8CxKbySNMgDy
nQ625IOk3LwPGU04KLguKc0R/XhtCfgjKWWlM6T+mOrAyBvvtkwIyvax9MYYaHZrHMOBDhpNVlDP
BRBSGAehzM+zDorx8pkDKAr5W87DGwjgdlFqcP0qh/05TwoJr6T+09jHn1rcDpyVrNQ+uY39CZgR
hk7NOJRGTiPFGmFoDsRCNnGlLor7WYwqoAOroQ6tKZvYaNL9mLcU8bEVhOc65/o2JlHJVf1aBhGs
521Ck8zkK7uGPd3zlEb4QfKSTsFJyGYVNeUDb57DM4zCO1TwFebJqDMN2thFGeGqyf7lb8XpIWVS
8ylG75H6UKjPbENoN1PWZozr2d5dynompj5WZ+u2U8BsZJOQRTh+MbWSI1YZNRGn4A+1WCe8kVI1
b+exOcOS3puTafaxbQPiUOqQX+rBLp9oAil6Rqc7pNEp6d7cwmMWy/DfRsYtvwbUSW88S651hJtN
XW2zbLmQ+QtjphcrmFPjw8mm3jMUUsdGFUedUMSTdna5OxtujAGULWAdLV6PkXcB/8clkRZJ/s1z
G87gHvyPoOyIXJU2WkKZzImOpdbdhj+FsIXCJ8SPhXnS1G0CVtecvh5QTDFYY5jGOP9fCpxS3det
C4JL0aSSxT6SW130JPJTDVx5wtxQeDwLa3tc0NQtTa0xU6S2oCqr9dv24a9UZSAnor2Uxhy8fB3w
ulVyKXrc+13HC9B1B6vRdFkD0yqavWUhywnjqLs7mEcTnKzCMjiG0bR7caBloi2vv3He/AuTHiIC
aDHLNceST2WkvODsiex7L7GGCZI0JmZmV/mgTh0DhRpaJXChTYCshkU+Eb9uRQuLoBBVSCl5bYyV
qy/M/yzqUqYceUlTppGm43DXK3rziHklV+ZGHSzFi7qcvg6VgDvVRtTiPZJ2++HER5j1vWFAEfH5
1p8LTJysliGLH78/7HNyZGhF1S1iSuBiKiMaxjCeVUFDQeKwh2iXL1kWCRh5fi6radvxTN8rEWef
hwxf+9Jgf3qxKIG6H4TyhA27VPFunNQpe5MxE7jffH72rVPeyWvKIyg2LuJNBmeyva+KFKUFGB0V
uJxJ3VALdtIikO5usMXK2h4NoPv/a6W0A/Rzvr9c40Im/7/BJky4ccqFsZUDA61/5G210Cfo3SLK
cHqgGNfXIOqo98tmD0p30SnguSMvAjRDrTb/E47hxI+FQ1EgcaBrI+Gl2VQj0u3SkyTTrZeTYIjr
Pu5JT9FIouboiuNXEiDKsYfdg4uQiuF6ifCg4Nscko+fwOPH5QrktMr71pB8K3MHa7ZqpgeO0oSc
GoQUxCOPzZ49WgVtV7fVrcRZ1R7m0vFJe5mY3jkA6g1DzHfka78A9OhnRrAUuVYOI3Qbikeyyhmp
fyre7zsVIfnlrcQWayXk/0TdC2qBuEGyuXKDIGOAsYcC6HyEgY8X9i+LNGbwMULorZ29X/sbzdOC
CW7ZZUgDMm6k9isPKHRHtxIlF45HSszLSDyC35anyT95QAb9R+X/ZiRPZJgKctzg7GGEHST0zYP5
XLF6zxogBSRRritI4SKJBPN3Ug0VWNGdE29RoLGibjKN8cBoROd1RMTaoD/vhmIqqPxdTILVfQZH
gl1XBCVw+tcK6s3grPKyIh0MrcoKl5Tn2ZKkS6xyHPMtCLU82EbRzP/4mxtGD+UTR6YEQBfjtMxC
7KEheL3CrpSWVp2lk8Mb4pXx7S9ljz62SyWwii77WOTXXy8Hy1fQH18I6CLVFmCKSCpZyURrMCtG
De6TbeqIcTR850dNaOAxQi8M9Zq3KaeOMYSdhLmJt8jkqjcT94f2yIg1Guo51iD3j+0vbXA78Dc4
j2DXuyyQroK56e8R8YmpeyWlEvRZpvQWN+PsnjOaMZkzx+0zryOS62BDoRMfI7gpkv8BKNuubhWo
7x+SHsmN8Ap/csEc3xQF0MXGpC7bMT8646RPmDhHiRkNSYlSQ5ADw8f0TeeRHqizmeBVGb/ENmW0
6SeOAyLTBxTCdh5RfijtrOwqQetlnUyKF5HtcigyxXacp/Fjhd3AgrgRS2nuHis9OcPJcWyfEKAW
uLmkSGn4KpDI58QgOxT1if0EbtJYAqb6rTWfUoVsLoAbNyKtrjxoUJpO8mMCxuvakhhXVS06phtT
I2XQptuACHsETMigYeq08a8Vn4PwXdOewnnpoy9mOz8LZUdfR5OzGGCYieWiDR5FFCP7zmCWrmKe
bRpUHtI3SEYPwlth+8gEnSh8nG2tMBjxG0jOlyIIUKhdNghG8X/o0qMHs9LfLIhoALF60yC/TUeK
UGdFQkD2AglEQzI0q8fUahofucWqo+bc52tHVt3Vtgm3jBuSmxmVgZ1SlWsPi1AuAIN9/SS4NFTg
k53o2yfAhPtsipNBcg1ehc5En146toI86Ig70chx2ohYaXMRvIXtLrBBcTgwCuAi318uQfsvD+Wz
RP/KXkb5k4Ijy2WLGT3PL8LfrfLezPlpQY99KE56UEHyDs89XjeG0wkwoioqrcg5Q0O1Bo5NAk46
rO+PIMGggeQjYHg2fcyXTWMuMPD0TjSnHz+ziDc8tgsBPyxCMBFVH2WGhfYdNzegJFT0G832KfqT
7hgp7YCGvvxLjvjDnPZXS/IvP1djcwXN7/nGMlkXpMXjzOwE2niDSNANMgviETfoKGo+nlMfwQKp
kPyyeNLX53dCHaiAZ8bHJ+1s3eeE6cvwwZDKfbOpCRGRQZ50zFSkMMUAFiB76udPmm9cNg7hgoRl
tziqpxLHo3RYYXayPY81NBR0vHuyO4n/qOU7pAt0Jk6gLLyVEp8Oh/PDeK9CE0IRgkbjtygAjQWQ
V7selTZFy7/SVe9q7T86rWuWlUW3S/E8zVURy7Y2YaRSkZD+uDF7JVw75OT9mVVpPRx/G5gjMOuu
8d5sXhLlmp6xUnvLYEw8KbkJIvmmwbUC6MKfhDfk8NS+1cbAItiiFs9V8NTyP0uLtxZEmKERqa+C
+xHN5WvLATWi5awJ2VGEagiCF+x4LpnLADnENIcEmY7tuwHnzd6J3zFPREUriEjRMr8V32AqzW0r
pXyf5Ru7lFSMGAJbv9LaDWir/bgFOucgNI6Txg/zKzYFNFjuZwzy5EgQT5m96usvZ/p7AgGAODMo
Tp6TnafIuwIMOLSqmTVrMTo2OiRpG5IhKTkspRRTqdQqeKGEbuQmyNDRVTBI0hLWvFg2yIOf/v3h
0ygAIUv7E5urgUeJXduj03os4788MbXuRlKvk38kXwSiFkFS9hOXqfw0geyrEVubKdXDHMn+ZuJH
Y0x25n45CTOeKby7mq/3zf9y9MypgDVJch+D7G39+Y6T96JoHCWT5NaTBzp6cHnUBwt269WObf5g
QOWVJfUdifRXo4upHT9W9sLPqBxE+z2hiOgCLOF+HpDcY8Xi2ZksT4w7r2lk9mMmeE+6Y89UHTWd
5XDi2zcMHlSmwmNFsgsxJDcYZLocv5+25umtb9lZBHkUHsuuVTcxEOhiNije76MufmMEgrsGojmP
7k0ScJ/90ct49uJieFsSQgqbLrL0+IuylIFOFvkl0m+enD7Fxd5H0VZVeS6MkzCRRLKT/lgKN0uA
Ea6Li7LA1AWuyCRcWZ/43BNhJUi76nxIsIk1zj+84dIFsmZYUR6s+LTxvsfDKDG195UIOP5eE6Cn
MZZwoJCIsF91lN2u9h/b2jVG4bXTUTTVgy5kXFJvc02pPtnqnOLGKCmnvFKdJStgq8dfRUjKfShK
yoRId8lP3WCl45dBpRdkF02t4YIHW1KxP9olXISpakS7CB36OuiY00+1r6c0RPU31sLe1np/U+z0
7L5M/Y0d/Rg47URnHM5wjsDfpPEZIN09GjIeuFPJl03vlYnY6zKcLCPz2LREsgWVRfKNKhe0l8qs
oT3c1xjWu9pOQ4v2iOArresCsixUlLdC7/ntyKCcvA44JMb49B2wdSKzltwlxUb4cn7R53W4pAxq
tOSna/j3ayOXj2SK6BVn10CJ+8+dWB+HwpKKFVjF96yXhuJKE6t3zV6hQq3tMU+2AXrISLxMW6Sy
kL9SxfmxbqwzvGYYiSS7qqvE2HFDWTu0RoXs016cPsWqMBg3hZ2h45NLwLck5H/QlRtqXgFMcr8L
bHpyYewX/wiMcU727zqZ00bUs3y6x28s1mQR0P1JgpmK5VQ3o53eXkt8r+ljcAaoQDYVFOjN/R2W
jVQZjCbbKM9U8o3dvTkrO1Sar30XlUrhGYiWbgJb47M3FTJYLQhmANwkFCmyUfPS0crkMCRgUnXx
xUNgx8hxwD+NqC+gMlAIMbKRSkLcoqx0Q19CDtDxBib9Fc6bFPVm2SPeGxswfqN1kWMsbZK2OUuu
0j7fMcfm+QxW97XKzgTpfuM9Op3WVmU5ckNJqxiurWPm/EOyQhaBDBJYRtqwlgsU9jGx2rVidrlV
5/zQSebHAys26HtfuyDT9Eo8UEPVKghHqY5Y14+zgPlTJXZdScH56mQU+fzDQR+p9w2QAXEmdNwl
FSyp0DfCcKGFy4cNSzol7RwVpDL+hb4m2rjKa6mfR9m/hvy9CXaxCQOg31vEa9oYqkk7H/yGzIsI
MdK3jAPh5EcWqqDClBoAm8xjXPapam/49mCtu+fFxV2NQCJEWJfFHHON75Jc7bAKwof947/BrGki
qHR/KR00VAKQ0pzc9po/6XuNfBu8iiW7N6ZHTnlAV/kcIiQV/rwCm83CacHzNg2cs8yip1wrgi1Q
NLubw6ZV55DbxAI3sSi6A8zcVKG+cw/T62KoKigPXYmifM3i2mo3XLOqDrB6ebNCLUhKzapqs9N8
kNcUDkHHzirhD2pr7lYpkml38S6hFe9taQGiJIbCrZp3XY4iG4WIa4G6JASe1TFwPlPSUnkVK5fF
8VWNZadrYdG184hE8R64zLli1uaLqgXoG1VszBb7tFjZb69y0aId+awnRos9oUrbH3k9JYcHUbYb
44AxbEjM6uWd0ZU7/PoQd9VEq/X66kkjtDR1EGfXroDppD0Kh4tfJNw7FZ9LkfzNgyfnhB/C715+
eNgvEpo5trNmbB3XmEr7JOnEmIN3tMdrMls3Zz8S13uFZ0Y2hY+iJjhG0qzEvPe70HzoQ1HRDeLw
TZSm04W8Tw06Lj7qth3Rnno3FFP4NhC9K5gairT+Tv1HGj2vvRGT+jm/i+1uX9q1Et6xFSTYqD6D
u3TR3soseDUNYGsC7xEfA6VGYAkiiWQRJBJHD7lgRrgzgEY2xe1WTIKfbCJ5DN9s+BmklpCnU25e
5PRRFRnpywrzz1zc9vvOBTC2XbMcHDT7yUNjYn8O5wHr5KkrnlP31FbUEwLBgWrhzusokoNNHoQ/
HJKMCvKlhqKUSerVW0Kz6wujSgZqISW+5aH1d8+CGTGI8yxnCKzEV5fMhe3HDUwIHgOjxCKOp6I5
iVBtUclTjeRxvMSROeOjfJxm6Jt2IDIxhEMXnJM36a+XkQmuXNPZDjqsjo0XoITunzPVp8pADMlz
JsrkCQxyZNTXIuBBoO8+0ZXuS81qEBzGIE84NZaR957DBilNpYNRbbexJpn2tXaPt0tS7+ErqHOt
Zdnsys8vESMiu3EZ9KejeDeBhaf8GL5GDth6ho1ZlinTjtWa5kOJgwdspQpQA9XybEfMAb35ED+d
oBGwvsHbZ3Ipo8tVBl7q3gAN0TZ0vYn2ZirqGDIaz+eANYcZoj3vQfTkEiu8MfWh5OfhdDbivvfh
2UN1GV1VFS+9RqP7D+5sXtOX/zXttCXdXo17cUOzqa2r+Cdug1KTU0Px7gDAIaC8nW2AdD/1XzOm
NY17zyhq0QgMOJfjsxDh4s+xYMu82dPyUGUBRZ4IgSnp6gNOPQqkmL6M6QINDLOiXRnHm3LSXHif
fmYHzMIKy8QZZoQMdCaInJ7DgU/b3ApaEBqUJmJBMaVenvgU0zJadGNa+ljLKpDOlCeGc/2AOK7k
zq/9pb6ZyRP8lmWf+chi7ovRToCaziaOft/6vhYDf2CRQnuIivkz0BdQR49Qwv2BNrcFO+rbU/+o
vSdpU+q/oKMWbaKeQYEuegLhefg8P23+7Xcv2HQDed88lZo9NscIdZyhuY6lBXtxPFoRz7fEQwdi
CnzEs8UqO539wBY2XpAJ8h1+yn8AItoDgcYCJcJpW6jheek3RA3/eQEQ27XovfSa5X0TpxIUUhjC
Qv4N6dH6HWHfWqY1c15J/kVyV1NCanKMKnicPZoNdlE0hEIcUeyXsUC1Mak82OT21XFrf0OT4c29
Dce8lmTYr5xX6XuyGpJY0ToGMc9cY0S0xLey66QIla6UFKFJEIvI5QSdBcDIkhN4HeILn1J2My1w
aQ1zQ16nz8EE1E0Xpo2tMreHmRfj/8Bg578+uDc/KfY93e45w50DwUB7cu8YFKAvqNfyufhy3ZV4
0bk3gBuE00VSSKy5XnqRL2OpdML7hBBWONKbwbbL82p7WgXsNqUvhRCVVlVId0eguozbkcHVN+/u
/sTE3LJ1FGZFX7oyHEhpXeitHvNj24MUcX5zSWst/QS92gMNGx9XFm6I+RXkL+OriKvqkHbEKhij
uFTY+auq9Tr6y9ax0S6zEYFpBQvFQEucKXOhoQ3ZCpiUlEC2uB7EpyHOLQAWrH4U3i3qCtfA3R1R
LnuDcdL11G6vH8RxDardUSqK71p/D1Xs8JmD5AUvi2HPMQGFG5xsWDtg+D7bGt1XaKeO/3X3qmF5
HBDxm0ch/iK32mzKgy2dOnzo2ft6wIQMdwHgRd1Ku8U3fjL1HrHdBD7Zq6Xt9jdls05aO6DUYu12
s8ybC1rPsCvUOJBXqD7H7oVgo3uv9M0vtWU3/sATfE/p+zbc1VETs/ufTQfkMyd14OnGmMqrzMB8
WY2fYxUS+S/wmu0YfSTYmUzO3CteYT1azX+q6hjjTdO0zDkbNavT7NwDGkTYww3W6NZ/+nbBYZtu
GUAFdIINHRjuZz50g3HS19jV5CnZwuSWTYXhQlNq/Wjwr+2XqgNm1grbifE4gtItGmEp+S31RSEt
aUkE3uXNKnbIsyEuJ7ACTB5gWE6o7F03Q15qAUUbjVT4EOO81FbIVdAdgTCEoG3czbB20POEkJJu
c6eaKWVQ+k14hN2zoDbSLR/uIvDCIrDwyAHjIKSmG4OkOMfVNcghr71bZKtopQ/+quq5jX8qBzZd
TNreHMvhfKtx+/JI9Wu51cCoHFP+lhZqhTbBPzOHyQ1Qynt0vY4eQ5gQas8M8LRoXOZkDRSGXMmQ
z2O8lr8+fv0+MOyUWzRdWs8jb92lpnB5oYYc+HIjM3B+aPN4oVekj8fjSKrKK7gsJtijP0d1h0lW
Jhe5PevqVjAT5YGgLPpbeRn335bBhlpdodKkKKQljh3YpRi73eF6G5KKuIycZf9tnDJo2y5ic7Hs
zA5UzLiZu/HFN63y26NGdkWQFlcAHJvGzHFaAm9O0MeiKaI6CxowPTAwUxlq1ywrU+YFpH2km3XX
EP8TI46AyDag9Q5VGbkCiuxhfZosLRf50wB626q+ZfVPGNqeJodycGfPXgB0vO4qrzzGneSAxVwF
UYZXe7ph62Ahj4ayJrU91NSFVbcxqAX56z3h18LrdTVg0hW6oiWwAPvB90aybRaMCeEvlI8zC/l7
WnNGoyyTL2hRtx08H6KQWnf3bW2yWGi/kpzaPkFH+o8y6M1dgV2Ye2IzZ0eVCwlDFNw5SJRBkHlt
yiBt9ErMkamFef6YApdFrDZIETeRxVP1G3836reB8YcEpjkogON2rLNs2HuryPQ7gRmMIfvozVAl
Ug+DHFdBGFY4gvbdDbFwSJSIxrxHBwQ0oBOb6HnVyYooHai+ahAyBD4eXjdsODMhl5bnOpQtePyG
X7ZYO0Cny3yF/z6xJ46SIOtGT9juRELFaNem1CMUAQ60foyjkLP06SiklDGsKIy1BaECoasP+por
nRBXAcylTywo6KVqjvyvyGf63PRglII7rsJEUq1Suo6Phmd1Xk7OYRKhpqJFwrD6wuSQfLDS0B+h
/OZ3GcyuDqxdelmkC/8qmYWuNsYkNLOQjUCi3y09CWjMj5dj5RikGhGjLuyNUxdMHga4MNk79oxf
ovwgPgeSCiG1NYUagvsvy1aEowqh3u48703gdBkxOUqlAPUwQRtAxgDLD5//jVjdCUmFoCv5hTpo
ihBW1gIQgrMNAvkEr5MTOgO66uo/vzU6iNRMhAZZ0feuaQlWWkLqPQAWZLucYBpgNNYQDlyEoymb
L7zgH7dewKef/WjtfBCQ4opbk+RJQcTV0gqoGvnB+bMM1XTg95Eutyozlopx06Ok+pQj+Tn4nff+
7P2LIqCjjdy+eW2bbxWsiiX57ciqz2c+cLcJChSiAa4bm4MkQaRvRZ/9BsGAEuk2D34mzKgAUim1
RNkVpb2Gnut2jH0W+VhadAw6YUFVT0R/B6qKfw6sjCpFSrLQ6TFb7a8KAvP3nOohXUvDGj2kPIY5
fHitDsynJCJBw4xSuSRWruA8qqn/a7UIgEjW8ZVe4ANGlx/7uL3ZQMDB4cI2UU+qSxddyYxq7tm/
owTr97v113grW4tMczED4c2yaqRC+sgGAe9RD2jPydATMmzFBD5VJxe5NJL7khnq3kXFlGiPfjsE
cymHm4+gZaH4N/tMFBqv5vW3Ssjq9Z0OcPmePSLhxPAN52t7guslHbYUsjJwBooyK1RDia+3FXfA
1rsiawyJE2Yg8jRTb/RFpldGMe6mKMdAZ2mu+S7IZI1Pg1fz1h5sHhWL0kxwnDr5FXqvoOj64r1s
NK1qEpZCAJZ/0uRYTI25Z/Z7Dxta11gsup38GpX4JVf9S/OCBaY+JXB2lz8+YlOzfSJ7dIG4PSae
7yWh3sKX9b0Jtxmuo7TKsUAChm6miqCNKZfjmxjnu7ek7VW1doO58/nxKCdkccEkoJ2Vpa7I4qM9
QIPjwxFi3HLfFwW16o5EtBAgPon/ttT4lI7F1wKGqgq5Bn/UlcaDwySDyo1QwG+bvPOYYzVDV6ZY
cneftKRdvg5txHL0X4uh46GkikoT185fsQjTZzsPAMHCl1n+WGi0uwt5tsl34P2rgE10o5XuwL4b
YLWGvF33INxGfcQcnFRwGXWrGzN3+VcH0cG7POtsLtnDtkfVgcQ10OCXwAycp35BE72qMiH2dkJV
sLMD9ddEQcd744eCNV76umBzghBdYqYS7l978r7plNGShJIJdQ1QxToXbmISFdQx9uh0ZhussQva
7HbENRPRYfEXUpegvY5UMKex9roSkAPc8JPXFt2w7IKAodNVy1SHzbTh5Z4UlN6AzOP9c8n+i4RF
JDabyE5Su4otmy4W0RUTHj1piy1sEc9AadeEd0GtMqwixNNWalrs4dgbV/O/8OL/pimdPF/dPwNp
/2LZDuCwAM62eZn70KczajgE9hoefuwAndjA9dxC7NEA0nneOJHobG8a9AqPdmpafby6WBaCKB1c
oS9JeLcJ/MwQ/MeSa8uQeyqROETEmEqkxeEPnGGQSDzOtyS70LXVPGtb6SsoFzj3Powgq23sFSqD
IT87TYiBs8x2kFeKk6xsAa8xXDuD8G4+orLq8178LXX822dEI+y8Ta9pFixc5irJWs8SahKmjjKJ
z8fDK2ntHPIgNnj7JVx5ZpK/IpeZqzXkeGsN8rztg3qhwBnWxAFtGQ5Lf0VCfvalJ47UBNCqxGza
LGAkbU2Djz7AYRGEw5GsmtN82rR/E4Py9pMrtHcKeXVSv3x6sSwUqeOlo22j0P4aYk1hfpZ5mUC+
XyQa8JB5k9nZ7JBsPAdyr0P3waOm/PmPf3cK+v+f15RKMDehtmDQ0bA+WKUGsd1MXowudkMAAmUw
G5ElrRTXJSveezYfHez/ZoZLsQSK1Tz66RDPu4trltZ1J/tJIAubXmUcsYuRRWQuSCG4YeECBCTh
sr3a7UqirVYZtAKwY7cdDEHeevLRlV0CNtgVd+HFOPjX1uuChKsOsG/L6/TXVTl58XEjP+hRL4Bn
nlvTkdrBC3YY6Ejdby7nyik5rrotFWvJrj3+dGaw+yJ3tGRmy1wVolZx9YUqVkSU4tWArnQ5NSuE
kUtMMeybuI5OaCT6qGpfu3S1C23lCegg3N3A0F/KLnky6UDVme2Pqe3g+zWi1K09MgG1OK19kTyx
xVtkI9LvY5jh7dDn4hp8DHNdot0Ys16L6nYYSY+FNoNW6W2HDqs2+9C0gwVpU/sYIHCqdn8KgMYv
K/UtPs0i8YZfyhxSwK2UxUIeF3nlVAU1mWhOP1ZmxaTKxvZ58PbSzE9UQseWGvpO5vhaDjRxmKRo
9jECD10ccx8kL5L3Vq+0XjBVqCWtb74M8DmYpPIkA2/XzxS56XHKqF5RO+cV6OcGMCnvAVe/brFc
G+2pCDx/weLkyTvIrVD46WlwdmW+HZlP9IVpQ+3JbSXcZvLvoCUo1n8I9Ca467a6cMryd5uIett0
c5i42w9G/AdxH6vnV2rWY9kWyOXZq4vcc3GkARE3YNISiWdodKiVK4pGOg8QUHByoIpMomaF5BCj
6U9dM1NdL3Nf3jib3ftSxfuXJknUQAjw5HrEUfxizCzjzeZcJX9dbBWyh5KWRHjKWKWZn5H7BZxj
PhYbI6ABLoj364LMYKThExrxLjQK6CJ57vD3OmwheXmWhGpSkaHQHglWOMRIo8n7IdYTaKv4Mjf/
5zOCFKb7rhOLr99zaiipqtSx/d3qwQ+R7Q4+alLoeZ4HeVQeihUbrQK7cRWZoE1+Vbgwwr9zyI81
kEFcgHh1snGHjCpiPgJT/nupkS784lRe62iyvCvEpSO4rMHZO1G1DmComvL7Lntdukfjr9UdCxKf
RGxBxq61++Ss67hky8lc0PTk1tnSda4amYoWaR0wLP5ZNeS9H3i4c0f0l0Ezx9hagE8mWgsNEIok
7n4pmFw2ciCs2d1U/lbsRKA/thdBo8waqD/Yr/N2M0Tz0IJgFE9/dd/7wF9z9I1CVcdO0xWSbGjR
WH5dwiz42d8efizOmEN8s+elNa4ltY5ereCVyL0opFmmS3tRBdMxtWtD459Ue9RGcuRirJPMiJKl
WyMULaGOeAfHesCHCd86QMS3MLAe4s0/UU9AD/3QqmgOKT8ttRhdWWQ0mXztM9uVQCKm58qS8uTT
YNFKybg+7UF7FG+V2AYh0FcDoge0mebCzDJjz02ngxHAXUalGIjYlGhvaegims3QrFIz4qAK+GKC
DJFgsENzvNhn67EViSJK49/paRGF/UmKfhntypuOMJDDd967atXOeAH7aatNs0H7PnZ5gGvQUd76
2rWZXFCF2qstPgcQj7gCe4tDfLSacvHifVFwoCDPM/r4C5qU6C8LPp1LlCbV+tThA3egENg+PK7h
QpIvPu67QsfQ4aa04zdKN4zIZVzhyymJyGPIUyAnTbks6hdtTYW+ChG685X69yVv7VK9uJuWZH3Y
46uKWl3fVWZgUml3w3h9Qy67eMmrVfk2+/JdgX8jRtPHL53JH53S0K5FPeklVY070BXlcjdtlNV2
RUfbs53Qq1eyWtTmkUSue/CH1B4yKJib2m91E4H8XxzPWy0PiL/9UyNGbCop7IIjShPr4MOnmMuU
N5M0W32Vj2UW7n7oH3nbLK2pqfhKjhJqSJawMv4mFYrFpeSF741SCsbOFsjeuAjpy3nufEU5m9EF
zId/fvmAF2/v/h3D+cYeh9elxvsrejwc+9bX074W1+ubd3FGewp82HbQCoRMVzFi08Ixzb7phj43
908X1UXaNCD4MG+SqvzaBVeRrs1LtBV+WnkIxTxynK28SxXIZzB8121Zslom0BJywu4MnR7qVelz
3SxHwYM+XeuXGnTKbYrIusQiE5tvqAC1jZmnG6p/zhjLnoPkpKfkRrFMOL7fqfg20b4R/I4+WzFY
Q4+rBUS6OCggbPEnKaOwuqK0V8vxclggDlHoDHIahJdDm/RUipxt/x0zu1opJi1JAOA5heqn7Yij
f67Vzqw3EwuN0Ln9GxVO3BJhQRtt8LDFcChvjwKz/ZH2aCfIzvlKy7SKGIytw9pe24DY6rXmbOLD
hNfAbS8OQBXvb1bmgfdqJ/PI5xWBBOjwdx4kj1P5jebQp0ZqA08ROZRVMV70/Cabis1exxlyJTKv
Q3pruROBJt7iuXP9Kkwcl1e1L6DAbTLpc3gom3ugtWWLAjuJgcd6OJbOW8CQ05VzzOpX4MrF/c1C
GrtFJeDyef7XoZwmmzKajgAC9sbHflXEzIb5Ap8va5DshFgL6rH9TsdJQx2Z99MCzu38QQ4Z5oOf
RzhRY6iuSbMab2zMkfxyILFfXux5yLj4hlZRWS9hMlGv8pqVRDWvmaGhEr+3N5igkJIJFH5VG3cN
N7A7TbB84XMz3droJlUZ9I4XtTrNTbbtwDLUaqSmqfES7/0z1aRFXnkGxLqEIEPL6F8tk8igDETC
5mSFaicH3QWmqal/ePxjRvC1K9khSQuwttlPjjzQabdRuMHaGiM660CEDjTGE9SxNPH3ybaKtXDP
hKGmfX2mFSHzYPxIg0gK/2Cly+4IIwx+xHCKOsX+1+C5wuSRFWIbJJ2FU6gzGukgfKyDplTKzAFq
5lA7HtNRVjDuzsqSo4xnW6+64cd+eWnPupSJ2ok4C/PCH9UmxEPgaIq7TwxOh7mPOlJ6osIJZrsu
xirq/+7cvF9ytuhrCSV46zXlcHA6n61uwlj9Vw9/Zn4dra9bs3UlJv13dlQ23F6T7MQppN4RoIYs
whybo7EIhOpK9tprL5EfHBvzIX0uc7g+wTOzGaUWiZqpnPqCFlx7D2ePPLMIoWpC9dsvrmjBsFOc
IHi7/XgrU0gr9QTjBlK7T529FIp53xJ4FNTX/OBtAe+2WYFG9l3jisUNW43+gJ3K+1jyO/wqqY6/
EaErAH0W6zI/AOIuzTc2OoSDCzrNktesJIvYvN5vs0bkh+IkdwXuLDGRlUjO0qZMOL1OWXksyDY/
vdizpMBTkkA8Oh13veCSEI2C3ObMpX5qwX4W34u3bltbniRPu22VRm3Q2CRrm/wbO0AdLvI++eFZ
dG9/k4S5Ol7aetaHrLAXgG2DPZh4pRCK+/WdUc2VWxuLdt1Y0Mu0DMD1hUHFEkuIDGE1GAd1iO56
uuNSFZZlIHUpxqJTmVC8bXAX63N7WifgDx+Sk9BNUSQUIUY/f6dbjE5VvqwQAunKbkJpZ9x7AHkG
IZ5NvkI2XiIcI+s848rHxj24Re8s2vt6Rz2ugkWKTaP1/tDnylFKCYPxGIsAOhN5EtQsVtbY6dR8
Le3iOfGuPWRge0lmSz8t7x2fZ4YuoLtpgwnGw5Lm3mjtsoLA1IA+KAhqWtPMLkBHUROrh85GnuEF
HWTFDk0Zp0df+XWQ9BfGxTe6uP0UE7RLuwhzTgfcjYsmk75Lq1SL1/UVDKbBH3JLxrzAHrhTrRnS
5t/8L4OG+yHVWxxYEpmbZZVZ9arKJu9QWHeVZVGCE4bcVsdvxn5P6Jb4Urg9XpM7+Te53jNhyDZQ
e7bneLNtL3Oe7Hi5FYFPaRtsJgHZ4RK6zCRqg+K8YtwH7zjYSI6f8qbwqs4+NULuEa0RtZsw17Oe
SErccvMyk0DbvYN9Z+SHErio+8pLq+q+B8iSideEJC0Mrik23Cfnu82Oxv+9ilcypq0rb5N6QnH7
LMyLavX4aDRatX2aaAyxr1LdkMB+JI4I4ezEQSibVFGHVMhULCKMQabKVRQB/7rnr9oEpC2Q7G3c
HOs/t2jgw3vcXSZu8nRk+L0QVqNTWI0nkvK9raSDzQLjhnEUKqON2Q+cdG3xpxvNq21lSV+K+ORh
kWeZTvj0JqHuFmUgdj9zDj2frGsJdXawiW2v95IhGBg+MxEqROTTrvKPb6C86dNy0bBE0U/g9leH
ZzksGWo1PfVfvefhZHNhN2TQo47kVqDFCfC3E17bZuFRix2n42GaNxIKVDxivKGVDnZTYg4AHcmH
Mh03ogX0kVOmo4g7/IfM75Q8kDNSonFr7GM9VvQ7UdzMyWedaMh+Q0ouh6eeyUSyGfK8dg39kyZU
mvFgAybhMbikfVPSxvDw6qDeg4mzBCmL9ch4ItuTBcOGRPRn+CdZYsOSkBHlMuymSLQQC9nu1+Ui
enZBKtbr2nXTp9OVePEfkY/KYZVks6eUTA5UmU+9Oj+ynhzlxwLMnNaS8vmTRY/dmn9mMUsYhePn
cLemVUMu68+z2wjK6g4bEmp2kfG4eRMaiz7/hto5U8akIBbdmNUXiRgqKioRXC791QZTOvrr/LaY
MyxsLzbSTFGb8k/8Q1BcfbUJmtT2zVcspQR+GsqbyctDSUqlsAlmt+b0zoIGm5toUI5Oy2zmJQrd
zukfTtDlPX+82RCE5akYhHXEhKwx+DWKjGGTw1fW9nA6cSchRG2Dd4QZa8XlS/RAb603tfTbn1ZN
zbuZEDxK1MBOh3V7MWh1mpIAOQQKRN0nI6KF/QOEFDdZ8CIGZZZZZOe5itshjdSQWwOsX4EqX2UT
thjufFBK+9Np39wlzQPxY0nZJ7VeTJRRu/bQ8qjcyzHFzRNuMQpc8Eo77AtRt88lAZuCNYaLv/Jm
H8KW9idW6xhw54Up/S90UT7EhI8bwNrnGg0BTCeKygvnZo5c8AHL+kL4GgU+Kj0Q+gZOG8N1ZV1D
ncdn0mwbOGXwARy4UvGkQk9oz6+vti+djbdo8TnkYwH4SatczBKMseFS3Nsa3/ARXiSCVoa8XLUx
lyY9ai3raxll5L2LcoiBvr2L+2GtZJpv5OpkDreg8FyH7Wpun5RgCLDjys54dCpo/fA6kui8RRlY
2ZjB0LqPfMbeqvXaayLQyY2tdtaFrfsKzTtcdEv+gTTnv1TcW63JPZ9AayqwNsU1Z9nW2sMJPUJc
P1ePwNhbrfR1rJLrVKUDjueNitITLEzi78P5l5LFc1s0Pm7v5SBqSajM4usacAyr7mjUJKrtf632
yxTtiHLUQFFoZGWJXJ2NhmitsYphx1I4gFvD3Lm4+iQngn21e5Kp7MBLve3DcRacby7+i4moy89C
m1c5Y5ibrH/UGUSOuy3zU8j7nV+xjxETyakYLAYVMXsc8sawvW7d96cXKnJCAdUy583eGM5Zul8D
Mn49malR/re5136TaytJ8kzIcI9lWo9pW5O8WXCCDU4gA5pJ3wK1nTxW8nf3ILVP/+K2skMgKp0d
9mEL0fr0MlZy2Ya9bjgUgKjflQ3JXyNFYkQOWfGpeqqdaLH6yXkWl7avnz5zltrq6uw+oBnU23JM
5LTey2f59cZCHLJmMuHQU3JyLgbDif6oQoBT73UJTJJOF59Q85lpy+EvKZon4sRnqlcmvgNhxtVx
8TYmP7fbBVlcBLtED03/JNn4hU/gdVaZKKXAToUmZt3tjEv0spspBMQ03XFGiWRdJ+bKyjGFlzY8
hZANE6+7B8gAKpt7a2knjUBJizgqIqOAkSGi10ouB/vA8szzLsicQkpAIAcrbYhdljiuMI0JSLmu
5f0fKwW36W+RW1qA1aHfbd7vaKOYBVv5BWUjRdC0YuEbMk0/Hnt6kPv85UuDTtJZxqwaGUFZXMbf
4LnRvwEkIW8M7oS/J/XxCkiUd7787ebrx2Z4qg6rwpISNcJQlGdspxa+4NY3WsI3amdZOWTEnO3z
j0t+xeP2goKrfbQyHOvpsdT+laG7xnefKWDiYINr/vQwlmL3PWmowGOGGe86xeaiz9mfzxDnLtvO
2fG0CMf+NdM3j+l07hs3BIdY4npNijXM05TsYWjp2ESWhXj6MopdRZ0KFD1u8JpiDCrFtQBxMwP0
l9EUwOyELPPpk6gd8XXollaFbBrV8cK0A/VOepuCPfiZOzuyv1BIasY3huF6zK8Bvdy5ZLKL/ptR
Es88QEphNZVrE8PGnzXXBkEfJvXjAzYEqmJSbNvfymerBDJGZm79T7YyT60fElf2Q63MHa0tP0oZ
33SigXJqJZRrXb1hlRxbatfv1SixUnZaqQzNWbwZs4CA0IWD3LZ9tCv+wTKD2SPt3FQux2GbCnQN
bSNQtswLmfRKRx5C7jC1tVK7NJ7xULV5lxx9n+KHua77N+FIXDnZVXONIT9oHeBzVEogIfmjwi75
NgCSaRyx9+/5DAEawxxYRZ2FCz84SN1xQ3UfN2gH4M9jql7Asa89eUOaz+dBNxVjibAMskGgahxx
exRHjb8BiX8p3bJSa3gbEBtsPesMc3hggXuF4nDflx52gZ/BKZ2dNiOpsAGDqDzU9NLq4vMbHMNH
6hrKaCrzeJYk43/sbibiZWXySdGIqomKdskXJ4UvPLfKxGjp0L55gxm5Pr5Bo6YLz/NFJJn9eZG2
LF7aIoQhwl6RjTav9/stug/tlcrsVn+FE5p3Txaxn7KLIpGxgV+Js5G5Gu1IjToGcoqVUuXb/Gg/
suzWIMEjyQeUQfjKgR9PsSLRT37m+Zb8nNNXiC+0oZFf0Abrerla+zQF7pQsa3mhRmLboWbfPF+3
jd6CNiLVxTcTY0FYXxEWWlY3d3nVnJB02qPz8gH2S+lL1JMv2K24S9CPZWy/CqI58t3VTym+NAHi
UzXtDiGxgzy+ccC7yMxCc9f3ZJux1R5Pxq7/XEcKPqTq21/7Lp4PN/+0EziudcqcPxnO5bz/akfr
aCYUVJ1r8+3X6AFsgMwISSEzqb8yFdZx3oqcdJEgo3qOH8xSpa87cWsZ142PiDN2Jp33aCq6GuSi
wiWgSRW9h/w4/E6CsQV0iSmzSuasun75pels9YH+jEScXnyZCzbctG99Ui98JgL3J8KNh3pCnO5c
iCQuTZePUhxEIVABL7A70+kOB6dgMvNyl+UjssOKosVni5KX7ULskuPgW1aw8to2du/FyNgsHYEg
7xJ2P63jV9g3X1/4M9PaoKYt4dbqoRH45F7OvGVKMb2tH3G9UtD59NDqgINwc5WIxcr0S05sN5Oq
tGNZ4tZ0Czq+u8jEggRRRPeRpXrPJBdJqL24PfgKnQtUeu+9EKgAzhoGOVMuJiouSU7glLhp1R8z
jC4K8SQHsPKfE+l4EioVRZ7Ng2sBo2rTYFFz2d6wQx0x3LmfQSLuA+kJrVQzFkVsGHkK8f4kH18O
DHSyhIfRAYIHcLaBiI+E8KsmyvZRVd1lOnumqKs/8NIp/oDOpVvbmCxV5BEBbJGuj7VmkDnhf+Gi
q4RH36NEKdzyOWKzMrDewyOeKgTLQJn4D+jYt/yMU0DyPzB5otpx6mozxz2zwL60jrFvsbuU/KHB
c53RScdAWJILSH42w0LYlqzHPpFmyW11vqAuJ3x3i+rf3lQ4OA6yEFSzE8fBD72V2cJXwh47dVND
J/k9sx2QofROPJqqQiED4GZTCaxjN/Yb26di8s7kAjMIc9p3Hcrd95NBaygqIManA1cY83fQFY0Y
kPmF7puNKRXAaUQQpDF0tt1AuqXoKEREoFD7T0nmlqyGEAUBvq06PcdSKHOOImipy6h4bwY6mKKe
4NWtUReubBZFTQYgDT3T9jnd3V7Csby7KReR5x5pkNXjlRcUhHGSP+dJgYkEKBQYMyv7p+AScxtY
x6k3clMNHNhQB0qI7JxlmRWfWtGuzbub4ju533GBWl2MNw+yz29Qa6wbmXtPKgubkTtq6rleWDTp
g5sYndM9MUgqw8Edi6oPt6YuF7Izd5NDPt4eoUxW5Gc1udR5qo/NRmhnpVUWNMZzR3oaEQQq50ph
jWFtZEbzWqGSy7TSMnsTrMi65PGPDsSK38uOkpyllFwrBfH1Wm2dp/GoIUD3EeHqYnHL2V2B7H+N
Fl3NJndWcw5tCrwR8gy90J5ivqUgvQsVc41wy457N+b/rrKSbwnu8JBcZLXsWehczLrMqo6w/ScE
+ukVuaD2LCVY7rNgWOuLezBrnoSsrPRd0elrLoPSkhxNP/1StPzocBfgNjPD5ZkiL+7j9QdYhmxx
iaBHtkqgJXtyZRq9FiAZjftogLSBCre3hrSrUEloM2+moBbrheygAoV1b5usXDADim+bqDqmKlRz
CPOAeuTiH9LDbY20VuhNsVd6FEK4Wg/K4d9s9IY0CXvLdmbvJ3K6pZCS9V2qc6EcAcLUeTP58y2i
QoUG57K5pakslmwwcv3E71gI98JHAb24tAwW7NSckKhZjsI/a6jgFTvZaDTyBPPLTgkYc8KgsMZ0
hLTEQ2D7sHZCszGh1VmfZjsGxl3We2ZvBbO+Rq4v32pzQlydjO95UMwzc8B1tUdnRXj7PrLFJxdk
ODiGk32m5YU2wW9FWXaKN50eOVRC8Rca04fC3mIXQceELlf0HIWexjjOzh1YspNy66a+LXipk7yB
Q4FB1gLjfC0Ec26/hIR17iT3KJiQeC+phHAxcNSyrhz7SWY8eS0zou9AIa/S7KUCihv33Mar15sq
5zDUmamJH6lhJd9NHYGGyw/EGeuxC85t2BXwvKPLNrkQcY2ritidZ6YJDQIIQOpjrPxBYAAQngJ/
Yaf8d66nyRK/fdw/jZ3pv8Gydwt+4bifD37wDXjsKrEONnAa/GnwnDQP+kN+8grBSg4pvhUdHoG2
XEf3/MouSamyMEqpkhumapYh/G29rmdHym9VWZgDC0SMeGzkuqO0kpnSEzDvPYsZx3oYHsrgCB+F
lZJ8+ptAZU6BWzbp8TTgB87mKP0ha9P4vamXxIaXGr6YN3iDdoeKrWn0MEBzXO618bpB2i0W7Gt9
u4tnooB7tqncQMcRVQjQ/g7RfgDJuI/rTsHMEoR1duC+et1IfIIzuLOVJsMCsUjgugRcnryGxkK9
308q3gzc/Ev9FRE+qj+mwEhXYKXEwFgpoyU7msOrbvtBvS3UREKbbyJjC+2FkNxFxkvbQoIzU6hK
g9MpZWyyglnvGQ6Vs6WWvvQHtqD9pTWTt0M2YVM4m8FAvvGTODD82sbc8qHJhEooHqd4gMFU3GCp
4eHKrMKCAAkP8U4y4zPbaPAna0fgHOayuu6h9nMjxy4SYEe/RzlCVrU3NMojfml5marymL9JmlqL
dzJezuah9e89XmpfDRma8Yr30k1NRqeqK0AZzcA30GnPiX1TZUWKyLK+OGj5eLx98FTZqP8VWe95
RShg5nZDzdIE+nnJnVTcssOBceQbMe7/QLZ0ACPvdiovSNMsqJbCc0v3AqM0PWhXujJsyvb7IPTY
7NjOXTJAYWgE5RxSF2jSh7yUViqYAZ16siwKA5Wx1mlyOZPA1zIuFCaO6oM+RLGan4FhV9zNGNGn
ssA45mna+lCZvD+Ap2S+LMKwebLFL47lPbqVgz+uAoTIXSFz/6gKUi6N4lWiMpmYmLXp4NfdC/Sd
8B6tGJmO9a/SQgCOb//WUk5S1t1194/P5HGMePJWw/byc1306svBOZyroKFYG0cTwM9q/aWxLegu
I0r01lAXa8J03mlBbvPmGv6GaDevwnNcfZM2tfR3cGPvTOd7/xIBCBdFbaPa7SsGbPBXD0df4rE4
K2HdfW3vyEDsgPE8u8v4xRb1jFpPHd3A/Sh37oDSdDOGn33mVQXRiylr42i3mdPAjClxm5I0tjbO
Y1QWI9y/cGMtWVZxLMadadawgZ8njTBA7N74+6l6EfD7CXyGVDco0NvWI9EKPgWpgbbavkj4ndJ2
JBXKHcyfi0Fc8C8yMRHbTgR/eA0Enb1c7VX4lBqvBN0lI6JBRRO5Dfn98Hr0N8wK5Wkjp0kJT4T2
E8renWPYsYbbhl9OWlvLhSCxJJrHUpfL5x8r07GxR3laQx7GcMLIQEbEH5bDh07NMmO5+kzDGBYl
Mhh7JMt6zWVuMl6lyM9wgJ3T9QXBr+51/Ml7VKn8WbLXGbWnzwswYxobEaLJRIGi5dDsunsHr/Lt
UYKLOb8H9SmvDTfiPoTHnlj498sgaqoBu3tYE4v6tgPPO0vGaE4SmJCnllbGhoVGyAHFewO6BD9L
ao9D8kA0EG1II/H5Y1P+bhe85N8A/iM30ak1jwfVKQI95ZGy5+i47G+ANsojjS6a7PCJom/Va85N
Ah5+rM6M0JTGFKtJhRMHqnmvbmEqc/ih2R8AJKHkz6goR18Su9FiNYfBQMBR7yNWD5hOO3TCAExF
3YYVYrfksJRxCrOC2/icj/ClziHatO8+O48DhslcPhlJ3L/rIkelzTyDOIPctp6ddscAzU4Qsluh
m0Wpu425Do1WLrHvMe2umb6sPW+TqJHqDI2eFu6PV1lDL+oKuiMkvPWePxnJJd+AYi79UnsW2i+1
/5gZnlU1iBEug/m15wXHD9SCWjh/T10qGiMEBtfNhKCWyQUJibQbUKXKzgdKvRY7+RIPp9ohCEoo
9+dtpqGLCT+8u9nadV0NPTt0L4c5dJRMsXOidlhz/rwNMprNdC1s6lguP4ULPfuf73DIX4V1VYo6
ILcylqpz+AhV6W47Ic1lJYYHmGEpxLasFnugo1ghch4ZA7IKDfNdDMEcV+sVmgza8BwSiiy1+H0r
PCXAE0z4Rmd2caHeWiaWmUta8OGIzQhwl2IgAXW7wmm+SRrNhyl7iln2uNvj/x+dwgTLdlpQLYGX
v5EgKQKmSWLUJK9th+8u1FbplWRdXj5y6EkW/c2O3LohN7JmpFATNTGLrR0sPdIqvu/3gvnxwlIg
iPg3uQX7w7Yej2SmSXwy2gZwcAIbX1ThYl8no80/Xa+RHLA+KFsVsXmLz6pWjtTWN4XYtcEjfbmB
HFI43o9bxvdzxt18bsO4K5LsN/5FGm4aX+6sQpsFAT0WlKQ5qrMRWWyFZ13KgAmNNwgVcG/wTSEM
2ddaevdMWOBqsh/owHud8m/ZRLQTVgRh0h8Mk5UMZbuQ5dGYjAio1ATkQ+Q6gdigu74V60k5tFor
8Mfk4Im2rSfgych3M7alIhFhTi2GUsnfFL5hRFsB9LFDVYrR72KSz5MnZTws61j6jRbc1C9Lzv2i
Zr7h/QeTv2SuzaL5wtE9mLSKYhH4yJ38SCL9cVh6mhRrE+KH6BCR/gT5gBRBQvb+jvbvg4UQbx1c
pk7Cz1PnkLHjMBqhZ4gGkve3W/vyjolYHxyI6EC/he6hvn7a454a9XJO3bEnjTTa19i+tt8ETo6f
FVdYUwhwV9uV5c7mzMy/0YLzZ8YMfHaOYWLRIj1D/073IWv7V0aIMbm9YIE/61c1+sX4xYplDVbD
auDkwIAK3aRDrvnU6u8wRnCVHv7/B9D9N2aRHCxXFJdJKiT5pOPXQLUnIFVFci8ezKJvLHR+PZ/e
4vYbFt6HlcILNA7tY1Py/1q0ZyjFn6VM5RJaq5J2QK1eG0/M0YuzzcOeMoIRRykoAgqr0zkSn6rB
HqDugW92W2FHBH1egn7g38E24qWFXMTLJ73l7eDnyjrMDHKmzWJyvqKkLzmVqHFoAOP16FqR9fjC
AbBdQDj/82EAQJWFr82/IgI9ylsclWVNZO9oqTECYyDwOQ0d8/9KfzK1FFmB3MpfHh5g0+j9ouw0
kmFmQzOT/TRdSRHY8UaqSYhCmfiSj2cBHZpunTFzga1esxUZCg5Jl8AexkD8SHCu7wI1bnc0jGxm
nyXEIqBWw/BmzLSC24ZtCTD+Q9UWx7tYy6DsNZj0EfM/YXQHUIpd1Zi4JQlwjm2mbDZH3l+308wd
svtpTvi8Ql5zBifMrZcdZ48x7bZPP2m8F3hA3Zc4tKcLTYYCcVWXwyuSM/WKhKntOmEkovUVwsZz
wC2reUa5ZR3CtuUO/BNJD93GLPqYce5RByvYjK5p5G+D/ONyFab9HEf44dImhF/BjUEzKo0QuRUB
ex57Z9gIlovOcKhtL3Idvx8dWYvwFSSMY9cjtX54IpHFURL0v401hUoxgS4MRfOnDUXzAD3vii/c
dWU/hPbdnJKh87oHSMHNDLnkmpLwKKd+qMgCgFRog5rzv3/5nv/TvlHtE6zn/tkYap+RbV1OCP4w
8PIP8Dxjn9DrhPeMZI6WQOudIaMpOECA1H9gKJ9p2rG4N1/ck8o/vZ3JdbIesWKoU5STqu8dn+Kk
+npXD+AQYxwUH7N54/ziGGImdQgATpw6aUJpLRLuOX3kT7ue+8VWr6GKErIUPv/HM1wW/oA1EebU
jA0MkJCkl3VJh9y4OXEFEM3qyMNuJsd+wvnXrhYJhjJgq5Zz31XLgF1XAZvqAB1nrnyzcwVe4JYl
ViBDU/eQ03JwLivvDdHtlrAS/VfZiktEAIBAghkD+nYtceRBHhbqR1Pctu/GeyyRs5pCpqrJarPd
i1hsGSi39Dadv724kG2YDwsb4pJhbea4ozZnecMSU8hgYEwOAxD2VaF59+ZkS7d2p9vllyPJb01k
Lf9O+AwWh8wEkk0tSEUrORie7xjMiu4+iBaB70JW9jzJsUCA2lzgSkp2Qf66kS8zBCa7twwcAQJK
Sn6gIL4mBD2aa+Dq2x69mXAUxqVSiZC08GAXEK08DjK8o+6j2KADb+wyrCgb6DqIfnKTAcqCw6CH
KYN9CzND2NzuehUXnAAs3ZN91UeIuIEDAIR7oQ2QZlwrnQPLCmMZ/M5yRgmO7EePmEc6ectUlMnp
GA28SEO5FQmOGLZuLM5fLV5NmUyIADafKeWAG04ILOC5Dha4fSuIJfcxfbTitif4DHoONh55e2nX
9ibq5vZb+S9yZ/jYdQxJAc63ep/cLyp5OBr5JsiEkroO4PeddjfNeAss7EOAq+P8vXI6Q47MZV2z
Ktwet+ikV5NTXgpziSEty5vs0Oa/XHrfux3s2FfDhMJ2e9mHDvlkpK504Bn94KDNDefURElv45E/
1AJuafXK3vZBe7YVbiMEHe949VhZXh8oWz47am74deux1+TU8k1x7GwCvPUWJgf63HXtdQ1u8gq9
pg0HwPSPTX+XL7JwmKNK5YhQyFD76rOvkQaYCm/bYNtx05XbIFQZR08UI6ExdamBSAkNWICGMB5g
1hjkykMy0yWx27fiw/StAk63TvbC1jPKuzaxBBUUbpkb9amjDAvorT4h/fIS6m035AZ3EPoChfa8
IueDmMVS9sUMR6xNnHNgT3UGuBhKqP0eXSPaxsyvPBrss81m3iLfo5poN0rGwxNPKShrxQSPPU18
Sq3poLIXPgv+/JCyNnWyXZIJWa+XNOghAn3ykzWCzr42nnVL4HFh4/B2s0rSOAzsOaVdi4MK22Gl
Ui53abpcg7MOJnwLy0msGqU7Mj/IKoSJk6GNjONidrgQ7qV/gQ/5jOZ59MzDC4EuNkbu5w0nHhGg
v+cwvvajdFvpKqYWve81nXdPOHhIvSN03kXX0SXGYkjwLs0wrq5CNPHEKJUtq65+N+Cc2Z3iTHbR
HorA2V6FkQiJatfE639tuOlYnNZ0/yadhFDbmmKpxB6MNxj3u2I+f35CZG0a1xRE5IW17jJ4PuVk
k0kWb5Cf4qAR+lVDFoCXvCLwKUAVO975T6wz5eafYdMhXMTNSVe3OyzhXncJCz9NgQyxw9h8xrAW
knJU+tGfftz+JpBLbegc4lCFE5136k8TJeP1/flN285clpMcd9wrXg0AJNEFomZ64kEcX/jnugw2
w/PX1B3zfwc3dujbkAGhnJiflY8UHr5y63Lw2wRb8BJyRX/17j9cNERPpc3Derxc+SQgOmAa3PmD
PbVjrv/ZJ0smKxMG/wcRhOb25N+50sjPVJiMzmuomfkeouRUF1AE8abKBWS+DVtao9YxOTNF5xNN
LShaWd07sdlM6AGgEkCGCgiXfLTwPALqxyRUe9lmHEPSYNBCG6xsXn78lb1pUmLkiU4WNkUTYPxC
g+3LEar6XzfoAn7Grid4Wd7hDEyWblBT5arVAAPAqj8himWY4TQusrKwt20DsCihUS7EzJUXqc6e
OF3XvpN5NQeEB1HlLzGAYhXv0B2Rna2dZh8vxhmgMXWXreokoOta7BUNnAUP/GXBQDzc2gC4a+bq
er8cY/a1V5fKlV1z+VFF4c09iJU+v7pzJcmsn40lhoF0iMLztjDuwqqPH7gVdnrjnUN3Xb+uXfnc
sgmZdA4KpTBw2/kFB7WS4N6dFSob3k1Wy/24EpBtBcnBlHLfOiw1gC68zaR2yiVGUFDg9C3zVEqN
cdhiP17U50p4DaX64oRIfJ7RWtOMnibtBKgEUi/t9rAg8AtwUSDCg7DXdbxl+FKbIbzS+2Tnh6X3
kCmnB2/ccCScbavW19T+luMY/GQ9hvJ8pCVOZBq1taihXPWL8IX9ycueyJLS2SY3YwHAti3Lr7Cw
Laky003AHlx4tNGx3y0S+ERnLvHnUD36ONCpz2724V6eG7ONPGCO9dbCxKejh1x0i9wmJqwEgjdj
BxB4yVwbOPc8gqqihDgo+8VBDiPHoGeoFJkS6vSqNYg+EWD1MzFsKqrujb7G2HIpCmhKh1R0YBao
ez5SCkZT5f+kqYInSCgr3saOJ5pjV1PXgUsKCxIiE8Afqu8CJRUvdfdNxgONfviW1qoaW3WgAhQ1
GgjJjoomhKQb3Fv6G0TRx8Un/9RJ0RsMpTOGY+5MM6RSC/dRy026v51r7edMNY1vjocbKxsSEVpj
oEoGQigJNiMJjy2rlKJBGJdKg4Y/NlK4zCjcEdyF/5BC2vh6EmzErCq3KR8t1ezWFQbeAsVvQEYP
yd//ww49692KQZ/DOxT+GqcGkPNA5oZatUJFc6iMXHLVQuOoJ754pSWEgLjk2VK/N/mLUlKe0XLl
RhijMTlOObpGDlLszViNlJaNDzU5LsknqS9yrt03Mca2K8bYZH60RoOJjwBqr2sED4W65XBulD/b
sQgQ2YhEc2Dvix/iMWtlK725WpMOEqo5DEmx8JHbt3ElhvCRFbebmCgNGzqCziwG3neTKJ0QCwNT
0o5aUWD9Q2qcR7qfigmoTVl77mQAZK/y/BGBTz098YVzo4bkRJHHwKhf5tMBeJV8rJlBQFyIqstV
UT9cIIwF/MQ4Et6j3Gy7x5YEkS0ZC7jARGoNZ5EmBNMIKtRb9hpj7AxPezu0jVLrRAQy6A5n1Tbs
qW2sT4pkKkrKQhdSTRh8OWnNolgPj7XG86obenfUQmosgDGzFAYcwJ3bk7nZhslMUEpODa2v7TYP
xwuVYtqG+IXrRjyOxUivlRgATeJpqGzOmBKCseWLWi+aVeYRk2VBgUuDcMbj7vr8NVILec1JcmBk
YNDkFEngjfCjLhDhEzmsmVA81pW2Y3GVylQg8DinPldiXeFWee5X4CIqU9GCySeSdwkgEfBH+79r
iTZMJbNf38695yKmSlIBalDGaM7Rz4z5gKg1IRyrRAc3oPj8G2+EzTrJPRejxqCg5iGz6zyIHHRd
8PtwaYwVlBD/OuFnbkiHkDczY2EdOUSmlsJYkuLFA2oygbPRhC0pcWPkbtrCF/63zqCMBi705sWP
Ol33zkVUDk8yps+aW6ph7hFKQhBbdzTW9iasIYl48Li33JrTMptzo87Q18NVSBB1EnmcHD/uVJVg
yCrkpAf2EBZQ+Wa9LLIeFoF6TccT6HAFC0ClcABivA3Y6086fYSZGZfnT82ebXNcZ89sDNproO90
RJGKeM0PBPUr4XoAq2EOEueY5H2yEwxjfJhSP5cUX/IxBHpycKxcHMq3qo2gUWTtjV6vT/ReFmp1
kk1iDuNC3Xo/OX86ZjqVfywUT3lmyJ75uZ7ogkDzLAHq8RcB0dGQ7kVKFUKs2rsTwkhonHd+s5FT
OM3pD5sYl+a0FaslxY0iwXub7BUSKDEzNcajAvw1sQDTLLQ1dSniWS79F2o0IfFy7tPl9AzO5tE8
fYt4yMQ/I4gRYRP0XT9cfwjFGxyV8CElqqM+91k2Kmc+a7ypOuA+1MJYZKAumT+mQAsamxCfRtBE
k2oLU4lwBrKYMeVs206aFpQQlPnJIYjBsvitvxYKA5rmh1cScaSy3GRsWnIX/moWOVKZ08Vx3cyW
Bsfl8VwP45SMW2hX5TzHNREas0fJ4THxAKylR7SYuzHzBXXmygjoOPigSg9a9PMTqdtSuAlqSTF7
/p0Fc5mej+AA5d7o5kkdijasy1LIjDMEEY9NwDu1EyNr0T53sGTVa7xhWkWqTGZuCfu4UNySWUy+
Z2K2HStQY5lNam2j03Jfgd/sp2+/jaFUXJ5Pgul52IkxrWuLgZ4D8kQYbvfg1eFaQo2LIfy7BgCl
bGzhh6LasHwDbedG3/cmpCU7cqI2yixVclhgC3g9kYwDDnuMvi7jVua5fRAOgX81Vksta4ipm1VK
9zi0FnOsrI5s00elekTasx3oaOB3wFEOVJxWSdInu1+7SDTcLc6PQ4bEns302dDeF9FrM+8WQiuK
cEGcRIa+94xeKLpYpE7bohAmK4fOWjJZHwCXwS3Yo6JYORWAT3+nxMGfrm9zKWQJRMMFb1cM7peV
pLttAX6/noZPvKFZdKL2Uc5cCySjora3bdpAu1I+MQ2rk8/rglhwLGlemEo5pXGuwRs39qg55sgE
JO8bs/uCW8ojh1V9R1v3uyhnd0RE771ZrKK+Vqs6DCUR3ZswHBsHp4TbFkVQuZSZcZH8lwuxCnwV
4hjuWCbGY7jQTb1elrAnShuX/OowX+1APu7eFmkUpvDvM1pO7FAVNyWXE7BeI9kVBb/wxmDpNRVD
SnR7GecSkpbLxBMlpNIzdHEoETOHGWNVq3xC0Kd4V/bM5wE5/VNd2RaQoIEMi3U+e0u0yW6+A4Yf
kcVrPOUmUyBT8nDPIhkSjdKf7f1P9mQnRMTcbjZPi1s/o4BScKVP8tujr+SCTVbvBm12qkDFMu/A
PMMi6LcT/lOz8o05jeyEDDTkb2V1FfNRK8b7zUbI0PoH+Z7HU7l+PePoPMxuFLr7/rwhvbPk99+0
v0cuP0odpeNUW5gx3whG8hNOIs+GG165r6Yh6/E+HoM5MLQmGonpp3mEMasqAPXeMUL9xEU752mN
ZStWuuT7DJ26NNiXGFLJRe8FMvIlwfplx16fuD44nWHbilaQ5aoqJxg9mgv5RlEA5WQ11x0yNge1
91ZUw+iHJ3DydpdOHkQD/CnuYNI8p84klVITChh5O0AVFVjgKqasz8juJVEL+PaZg2M1CYH+l3ob
w16DyUQ3LXpPS75Exmy5F/8AI51qej9pKbpvNP1MWRiMuaLC+Y5nw4w/nSTybX6PgyrbhREqj1YI
o/3nE+o2QpkZ9EWm2VwFw1kVRJ3g3zR9urgs6yI+oUKxtse60d/RlOlInAb8H7WHWxbY/qNKjrKY
ZQwpXCPBSPWjzrMIZMJYKGGl0tcFb+pNQzomgqCOx9eFpQYxx0e58HUbtLzxtQPsTafSueBXtTER
Iq2f/K75YX684obiA9yDJF3befYX0rcIOLKlw1NmKwVvB5Es5FvXRSkInn7Mp/p0aHRcMqJt/TqW
Nb4ooulyKuLI67dJr5QROMFhiX/T/x9s+CHGtpRS/c9LKNQs3HVMylXzKk8WMMdnvr6RO1g5jvuV
5UudQ1/5konxWWMqcicQLtO9suxQlJbV3whuZWknGPzR/7nlqG0Mq39rBPGtEcrhoJVHz1kz7aX0
6M21aY+jYkqjpCDj7pfEEbi+/UIZ3Znao0h6v9wZmZ/RXIilXPVpmJoV6ikVn8s9uaxvnFypYFcE
jWVhap8irN8qECWUGhCmhsXwMDqW+fdCtI93VkjisXByuq5IlwDI9GrXKqn5WpXxMpMGLG/Fjrp4
a6/b+vH8m4AJiuO1Fs+sdrNBCsxqq0tgW9b2LXemo+Ce+1t7e5IEAyKzkja1haW+HEl7J7jA+JIj
W67QohI6gb7G1JOkO+aOSKb4g2ycG0DE1I9jMaanj03kKvVWWIUB63aXS5FpGfZfwiXoro1XyHRH
hjFCHoW6IvYgkoqxqzr2DwIkiaakVCLt6mXJvLw/Zdl+Y6diXnaUkkLAW5NcaIJUjt1RoNWwlaBb
vFjxe+0x1u04YB8L7/OzRwOQd6FoY4TeQIBNRA730b6Y0h+fIWLILmA9+GlysILVF/nvAenDP1Nc
S34gOg1Lflrib3HqicGgEKZwaFQ5bKZwYfHfPyHdYcIkc/7RxiKgXrfe+g4Nt/Ry8u0p2CNeOa8z
ivM9bEgiIfEFQybFR1WowUkHJIs2cJvQx6uZbv5ISJfPHoaG09qY3XoqSWT885Jkrk3J1VKu5RL9
4D//ihV26VOckKIK8qxBgvtMN5HkHmbyiX2apKkLhvo8/EXZKZZiCYyYxTLsZS8NbGGWQF0YBrLQ
+0NvhYNR2LedL/Xv7FDKWtjJa1W3/D7F4UbZu12uwHaFm2tINE8wsDn/9ERbY6dJNVUdGbKa3GE0
qPUPQP5mwQImH+YFomej0/KItJTEhTRMMrb7/x4o1u4VCicYTgwB/XnrNtli3VruFk/BZS7Kfcp2
Ate2yucs9PXsFCbx5R0lHfK8zd3kVbbfq1ejmPPSMoZlY9RcYg6an2sT3dCcWanFg2fOG9+GUT17
jleV7lIK9vMRlZYBsjGORvoZkXJ0vd7+a1srGXERqWCBFq1rhhOkDXL8ibO62QqY1YQDDhTUeEV/
LahIx9DBU1gmh09UywUehncJoviUCZ2S3yn2dFJ/XGhqz3vKp7V12C530hLUANP5TkNdck4vhDRB
1pQa+yBW26iCSgY2l4Ta2w/nZGDHwbUGp+6PJQt+/Ct36TgCzKdxJHRos+GY2Y8AY6AT1B1Ua0di
7VUy2o1xb8pwquDYTbTkFUFG1c/+og7sDri6hB1XEWeDHtCRidna5vRWuTqAUNwKcxstV8BwHRat
qjHF/PH+0Dc2MtAZR05ABSmWwNnecmBl/y8OwWWAOxpjVM4gxTes9snYdweKranw6ArzDqX2mwTO
o1Codo+49YQnumHkkTf/TSmvHzxEKP7Ewy7QEaMVKY2uymb+C3cUAd7WthT1CpMz3Od1kTznddEG
exdo5D8wmO8X6U3CwJDFBApn8Vg4ujvq2alKYE7xA232xLzqlhIfZTH7xrdCfDVcPsnJi7HgN6QM
YXJZVMQSY+ruSdNbbI0BY39xYg1Bwst30sJL1OhmC3cpKqRZ+4lpZjfbAzCHkzjeXcsKSAxnbOlD
lxfnh/SqbXUdOUvH0eZKXvg4c2ICjCeBh2cBE6WDk8GZIfnByAfRAgvB7YO8yg/lIjKvN/7jhAjG
npXnsEAfp3by3oicYESVGeg8r+XvhROsJBqqAqUsQ1vZWw+TZ++ysTjoJ2Ht1EuCaiQwnSQnD//l
DkUOdcN1XspZCChy1JauJhtr7bzSF0E4ezsR4SGywn83ZIHoLAuu5euLqhODMXfa4c7p3LF1wJhq
WCEewwg7yfE3/5uYwnZwQELIbGrd86GOYLp7cxVViE673FIUdKhRlzjqrMvT0hySNdmLlHfQjeMH
cc707CCIqkoskOycb/qNnMayR69Bb6lriJzxD+UiK/BWdvCoDKzv7FCRw03jXoK9QkYd83os/AuH
DAydcOLuXtNgtSUUBiolPpkYtgW5SE0KcWi+lhLhpguyHwLqyEve15eLmIGG0ld9VNmt8qovZ9Ot
ha0jYGkBj+2lYqnzXp6TduMqiTKrz9khcFfxpuoBUmuIrs0PvyDNbGmN8wk61eSK5LRfg8dduxHM
+0ErFTSudbMf1YIKKpfOYmEt/ys1m67fZsXoY16GMq+RK7CjIp2WgKi5eLeOxciliOit20e7c1Bv
3/khI/qLhP0hztwk2ZIwkJWrT+YR43AyHLTJKoE1MzNzeMas51isqZms8Gxj23ZAGhOtwivWtfxp
kB9fBj6gsvm/3FuHEhs3WDaXGgaoLDZeMZ9fKQXBHFtLValVQaa7Pzf7H+Ns+W6dexu+PPfwGUD8
CALFvw2PGIchwLyxOxbv/2HF0NAhV4rzOdX/kVMvCf+mFFwtnSrSlOLO332C9qnrWNAIVhPrsUiQ
etOnr4aMlpev/pJ5Pp2jbTG8Col+Uy6NzhkjrZdfJnEaK9gic3+qV1sAaM1T5lChJQzI6bVeLpPQ
5ezd830Ahb7mjx+UQtFFuR4wpzxfz63RZoooejTil9q94ZKw7sZUxgM2ZhfoboadlQRIj0LMYNyD
kPGhDB96H86gjrL7H133xac2HsZUDaJRzZzgqKr8DTpghUsiam5GyZZfL5AS904qUoU7aAXBLUMQ
B3Xygt+tEks/3w22rZTUcD2vik/uWMhETJbPnwpnUZhcAkhd1nTGz5l2airPVjBQ6EmfWugRggy8
3Sc69GDOm3+FT1MfDU2MObpJ8BEqC5qGgXjDy8mgbfTKXTPw1YWAlvZmX6LbWioI/nHVqpBEI/fV
BLsBD3BOda0QNAXHk3vDqllA0t4IvzpDAlzJy/ateZubVd9oGFnu2+3xeSkijMzg7KUTXHmeglG6
8+v94F79mWMffJXjZ1lVmwhEdsBNyNVg/7nT52AWTz6kvwQgs16Ei/qX2zBf3nRajj9HzgbEmpQw
zrxstLnSDogFDRnUwatqyqvy2oGVNwmmLUTxFin/Q1FcApUEjEitZ/Kmotr/FS+XuOWkop4C5XbK
+XDweYK6d+MRo3Yuiv3sjFEDKiE02yqJHnELQrVI7aV4cJBPXKRImJntfevqHjfPSC8uBB8bOpmW
fUwxX1EyRnsqNMwmHiVWAN5GojXZjwlIgQjGYBkqwijun6uS+/Ii41jS7DjcXQzQ5iWsFyqfa8ZV
ojiJ7ykYLRLzE9CfsKBnB1SD/EhimVVMbH0shOO2QwoijMDBiOS/TfrvmcwCxY9r9e6517KsxMYX
eTRrdhGo6xuSgCnWleISIrOJr1QQnsHhaCX+vq3jwHfe5HRQJRr0C67Hsezel1uD+QdnnHv+gufV
bDJCFYtpOQ46iUiew7pjqUzaXW6VuHkEc+i7vDyUeqi7Um5+ZXwIc88Ut5PdBbkyJxWd+se6Xbu2
gG8z1/bazW049ENsw2YwJbeMR8UeoI2h8hsPBQ1pnP8kBbOle/ZG9EYR/riSnt83D0vYKdE36G49
pEtI2WXnuzztx02tLeSttUQ7qEcGSu94kwlqkkHDM9Cx4IU5SInfNLPuB/XONCMZDANM8ReuD5e4
wXMYo9DXMMFD2X/GJTLg4mtb0KGMMJqS+yJGbImIE0MXjE/BVb8Sz7Vp2k92vrDf/0Sqg1i4TN9w
WIU0hfzQeSU+n9aQhX/UHf+hSmDBYVWwg8u1aA61VoSHA1HZdCuMhrVPGOvPYIRUt3AqkfXGHGuD
4oB5resCGNkr+pKSHe783O1sEyk9c2QylvRLHRDriC8IU6ziHjYKhpC/bVHwBOUbSa2hEstVrd+X
r00I+qS0yffSGkswIgnn1+kJWTsnZo2sTNk8xuonque7veEBK5dzocQjZXKnrixmkirvyeVFbUF/
kCLCgp8qG2Mc6Rk3vD3R9k8PM8ES2jlfvPWGL5+t1JF4Stk78zbkF7UO/NjMmbK/jcUeei76imtC
daQYc8+7jB/CYblHlo6jW4of40JKRWEQWmhv9QL9aVfRBcthUwkKChqsS/EP+ZhptYYXo0VOPppS
NwMe7tEhIKadgLNH4PQZoDbF0pro9jrueemgRnHz3SR/ODx/kQuwv8vlwNjfCOeJ16pS0WEw6Ll2
xK/Zld7E0E72HKuddLVY/6hxoFU6nVKc7NEpvuOuEwAil6Vas0lkf/NbVGgisBVBYmM7C1qYE30r
gVLKStRKk1pVHAOSPwfmUAjbA8FYG+Uc0EqfBioz4kBmtBJdL9crq+7qOjkNElOHxepZKX+TPzIh
4LeC7xZ0tdvvG4M8vEQhxA1WuAW5jNvgdRMyhE2UsVMTVbwauexKouJp0tZSHocXtp421heHBiZn
KzfxpYNRtGi7qj9Wxmj4zxKi9U6jAsCu4miTSsMcWBL6yWqvHDjtnEvFLDnZDsrhT9qlG+9/GKXe
1M27tQoPZaGupxCfolbnPFHx8inc4SkHzpSzhJQPxJ4Mj4Lt8Fsc/kO/OIZZxDin/aJfNmTeKZ7Y
n5z+I6tq2DzXDFDzRhLkJL6RdqgtfZ3FlhGB6tBe9ZqN9oTXWg5gnY05DRRsz9UnpyN40S5S4SwI
xP/PqCApyt8NcWJZ9/Az0MTLl39bBUR+URROVV57gqtlDcKewx2HzFzItVmAt2sMBeHzIAnK7ioo
la2wNCGbwPXoDMdXqwm2ik9Umw17i+Pv5w0tb6e9k0R8vQkAlVsFWlPQFV7JDKtuLoQ4oU+4na6z
N/MQlRxlCBWG7r5i7kkCy6izWnmFQLYnx2AjC8pkeelOrwKV1WtTekI3s4XKmQLFgnK79+WrjxV6
qSVzdXNMiXKe6uOpO/guTK10nmL9n73oKQeaKtpdB2+9AYGCJJ0qTfQU4LQr27FO06DW+DHCORpf
TlH5jmR1fHRNwKiIGcqrBhBT6XPY9M2O9a59iox8t5v/LyOv/5v8PSGYm49JR1qN8JtNdY5ZkRvT
JP4ln4e/a5jN9VF2DMlvfK281OR5/ZM/DhVANCaOqLSkY1WDj1k7EifJseAJKcOvj+sQ3fH+rQEQ
Oc0ZGHo7sxhKr2ZHn9Rp3hbFeT33iGsjSEyj1ZGe9X5sOegcky6q/yG0ug3HoeklqYs6MDAzK5Kw
Dmklvf/8sm4YokjMxNXUq85IB0hXXMUNiX/eRVwN5FUodbJfBMWV90ESwTfdVPq6savdOKVJHqPy
9KEJT7UOCLqltIPZmItDfD3Dwm4wGFO9H6LHxMRYYN5kE+LGjDr/5D55kQEnj/CgZZtUBm/wcwsd
is1P8gtovaq9DT1egI9TnLAI9lzibmacIVr4znFCAeWQmXaL3NsF2LAw9zY15e+YKdnYVDFDZe8D
ZLSkhXnGC9shWA+eTqIk4fAfJDwNl/bQMRDPJXeFxTr2nHHAHlSZY7CLbeyE9XJvgNINeQySeU/g
REsUemRJIFviY+hRe/uox33+YlTwHounEe3n5sNyDYb3YwYt2qq+4+UJcZyD8aSdX1nLiRXVkrr3
dQL9g8KMOhS8BS2g22YE+7H5YFzagQ1n8ouihQU1YY94+Ie4z0hs/yWqHTBkhz8EjUUt+hzwrWZu
wk9jwQpEBLD5fRZnrw4od4r+d26kFA5vGr2AHAz5uar7BZG4CuKYNro+R9b0UwvMNyG33oX1LypU
bUiTwH+Y2j5wsTPEpmfTcvlGlQ08MjQ1AeD+CAX3pV5YL075kgnzg9l819xnu7Qea605DjtVGSEv
moGrbQOO45w2PCxWiA+AAk55JVbyleZhUzgt4DgsIWhaBGM93Z8+sT6HV9ER43vjFA7a877GQAHk
9OsjuKkezXsJwfoe97LnOFlBgQtz9xnCxju37Ti0G9vevdEDLOu3rOPq2ywzuA+TrA0G3KE8ugVS
hcE2NvKSPO6C/PkRb5cPQb4OHrkiUB/9h7Rk6S2JC2RN1mEeKOL7OD1zCygvreDy7WI69/8mPeif
JsBDf5uDA3JXpK86IlTalcm3YRRDfXkS4h5a549KKwZVZZpfW51ouISPwAglhlz/DQh5hSuUDQBe
x8hDtQFQf3C7mH/mueZifsPO/cNdGz0rMQQF3kjvJuu5N6qea/DTBfNY0qeqIjICDU2qFct9LES/
9v2VCdPwzDCEQA4rgH7Lk0bzi9Rl0wB4fQot4COsjN520DIQrf07tIGqQTftxgrioh+dS8gP8ygG
RFh+VdxMb8mhWRG2399fQ1EnB12LoJCBjYeC9cFFXu/0x+kzTZZy8hEFhDyUHGBmeSUOkYKjYxFp
58VO9eX9Fe7n1hrCSwTZ+FVyBvAWHs5pCo0JYQ9bpantjQTbTvTirExLeS59ej7Yyctg75SJ4UDr
2kpLjqSQEXTlFKYMgPNL3uY2C0F6lL5VMFho5Pzw6bWhfa0Nw6ZAFG6SW/Tmg9J3VECWG3+eNRq3
AXAi+wfRJfTMMkTLfcQrNwkqdBCeJxGNquOQuQUtCCc/UX4x4SCFNb77o/EvIhew4BoD5eQ+BJqJ
TH/0MXMxEdmjmWVw2u6fg9AbBne0bhBq+DpigYjlsUVw3yBIefisSoQganFD3KZoAM2aGZbRGRO3
mko+akGgrBqP+vuoFN0UuVCpftG9JqU/nN4E5LL4C/HRQQNyf+IVKjFdRN1Oo4Sbj6GBRQ3cbvB2
fqBdgDf3G5K5rasV8oULGb9XNOR/ngApMw+riNHMufoz1ItFveRYsBqjHSCqdd2tMWpxfZz9yzNx
j98bBQX2cwul9RQSDByaIlGkfymkYkliO7cNeXMCDImxdMij0ZN1Oj0yUP5EnG12Mua0Kzbej+V1
RXUGJDMZqt2dSIU6jvQ7SH3UnzyreOp5/G8/GpAaq5F8s1uZDG7oMrwt/Mpd3HMVb0iQg300D1mp
LCsYq/7ubrq/DDNNC8Ui1J29gikfvDQia7vFKAcWvJ1C53ImD2m4I1Jm8bkemzUHptTUEJ0mQfeF
VUIQwNnEqbcRhkeGR64rP9xRdr2BGBH4vWRhtanIf2fOFLsZUgfFpTsVSLLu6gY10DkP+qDAf+X0
HhA31xhek/d3e/5TcJeXimcvVuPom9/57jvb/roS05gcte5/RDWY532CYf6+GPbkNLUW/EwqJ1OC
kNNKKSOuk1iCM+dT/fl1pud4K8OTyIAGX3x5HutFVbk4YqWe6sKe9g1rBQAaLKacV3cJ3aDLX1QD
TBc09OcqLz/RMsS9MQQ+pBJcPPqdX3N4rQt1NFDD+ufy3M5urZgmG5HgP7wbp4afqsXGQJGznAl9
olX7Nivoqv5oX33I8KmJUXYkehwd4iLzOj2tgFuX++cyFVerOpoBeEhycj0xoFpAlx6W9XK8E2BT
S1w5DZx2W41pZ5TPaliVP+4yZRFhW4T3sO7WQs8tXM/L9FNbODUOXsbCLLOQ4acM3DUNP5whtDUR
1as9td/BRQD3x4mnmlu8M5twE5qkpZFpOUFt6FbYK1ePJIpqStlJxpl3bsYpuJobxyULLqH+dDZG
Roi7A97no6qszmzq+qAlP+x2GHhpnuDgwnKyAIYRiBUdUkk8bHnRZfZCy9aaqgR27KH8CZcFE5XA
8po8yfajGjqOVCj2pcr5OtyAAsH0gNu7FUxzKb3SEDSo/lhm0h4H8OonkhQChn8i+ZNkH/ECE5XJ
RsL6yLPB4jG7QyKfTlzYFYbTGD5GAMWU27ezR54gEvD/HxgaHr2UuP4MrpAVnUcOmXQM6L1CIK7C
+KtwdH3oJI+q2fVTQZn9nFC5rIOcCHdexLlsbA7tUyX2SmPsf+wsiFh1PnonrpagAvQWlLlqksBz
LyBEm05dSV1+8b+BYehXUpsmGtuOrSWoqKg+9ft7XaefsMFL5AxvDD9/Dam2DXAib50JLHZqky0F
7sDz36Jj9XZHruxxZj6TKWdQ0HKpeVcRj4zQfA/3I8+L58GrlnzdvJfuinUv852DDC82L4JvvyrK
uaA5WpyN9VA94OT1Oh0IpjieYLNKjwgp+lvqZGVVsU5pH2Ya3GZVNL3/Lljk368SKr+zzKs7EKUT
q0pEs60cYksofx3HaFZaSnBnEY55hdzTGDihu2jcSyV1NH4YINlu5doXNgd5qGtnFo72UDqrJKWM
sKYXCVqXOubYt53YNkXbJ2yl/mLcwBAhBez8VZnxrxMAXsbjHS6FNVw4y21IRmMUxovcbjELl8jb
wByTcJyhyeFEAaMxKDP5sHGidC/PX601FJfuxvcwfpH8foQxCDX9dUOq5bObMIFgEJuZpQF1uKim
x8x0UsWjIArUMNW+78rhh0SXMb2qiVMMev7DzsFprzEMZ6kj1L5E7wHjXuUjbvl+8+gVF2mb4hKV
bSB4HUOPeng0xe5GRspIIzOZqnDL+rpUS3MFvCnX4PfHU7BfbKtAjsTKQdKIdm22u+oq/Oj+85TN
FPv2PanasWbNsT7USKabqw3ekaUwCyWoHS4aqE+3EBsXMwxtDsyF6ZOAe3KuSEBjz/tzc5ulFBh2
cmuSTMqF1B4zUspUhjUhEep4B854MNHH2GWbXn0T1C8YYtVL8/aRFG9e9dSUQhg/EuzWW/vYYPmx
QsuYOG1Wjh2gwXgMHKxwLl8+EC2XMOaxaKgql2m8ad8ZgdKmA4jlMr8TohpmbyEsJFxdiVugr+lV
KJ12pq0x7bwIqAiTVQXIZxeeeepE/KqMatHOVM+kALd8XtuNp0lOt0nPe5H7MfEosLyUR+5V2y20
MW1TCMLjponnDMz6DgEn5vZS2R06OTeasNOjpMqXd8wnqUELb85tOELJkOpzr6xz6W0P4jYOjzR1
+YADq4a0LcP5IIHgjSpdLTM7vjrWiaF0ZQEMD0IXONam7m7t64IcZsZoBi/DkhCaAm12qUVGUMwO
eshWLzkOknNXO2t/PvfNvDPypFGdA3KQIBfeqcO5rFGyQBtYrKTQfMenIXfoI31h2W4Jqga+Q4jt
Jyg6dwL7sES6L/uYBIFxU5MKQFy0Pk6kOQufi7wWsQ0kh7DNu3uBy+QdfZTR4Rp4SmKZnUNTPx/w
OnaWFQuQK6ZOlmlZTbGG4Ld/Fck6mp631/N9V3dV2zFzLw0k2lRBaUZ7Ig7EzFNdy0mSWBkX4f/r
ThUCgTaM2195Ra5rBc+Lef/j1VJY1nluD2u86018ON8fYqKgMSe5ZykCZpH3f91DwgV/VwasLglL
2SaD0hEUnuIbFKy0iFhi2Pl/zTItDWhu7YJ5q18ZWEe/KybjhRB8IX0m7hTV3LZGOskqkC9dLNNl
uYd44hrE6tkOvybfh5wfg0jLq6qgyMvWr76i6IWIjx2JnwbRJEa58Mq0BaeoiyDp6zQumEBQjTBP
y8CduzNPmrmgxXfjy6CoWSlclMwc3sG/QF8JVPozds4Z0QhT1R/l1U5NcZMsyTLMZiA2uiOFrdJE
9z1MyHiBbYlT4k8FYjgX+AxbxlfiEg3GfUa9Lm6oBHmhH7/OAaK95A8iiNJj+v4u/OW5Z5d/GVuo
EV0jr90BTzCy2fXvXc+3JPWfWCRtk4kVknwVq/fhKFegVXceXBgBg2dV/m5zkQR6uK9xkvMGWJaF
vWQoK6jUScgtd1adIIfc0sxFlGbjZBanu/BRGdDdmoZh1TpUulq5Tuc3XR4OyTeBPcjODMhKBYEx
IyzJOi74JeXdTMsIEd7pj4jRr0I3WpIL1EDUIKOUWrcEbVNHVkXJX4GQdVxxYBgSjMdjFaTMdlhV
hwPxG3b2y6RgysA8tpCJ8h1kMAFn54fu//z3CEsRUZanIr0vWXrJqvx72Vx7ybK50I20on5tNK4h
IQNyQj+ToR1V+xbna3hx0xY4ICSNsPCn75nPX4HFS4pG+SvuWvx76CGi8ij6AtJYEA1BQESIUwZJ
cnwETpHUY9SZhVMz+si6v0CtVfFkX1gxkuauW9vEVbsPzSO8Ny0sLNLDFcIjvP03oqsBLb2cKbo+
3F+3hTSfp1OPn/8HELuoxJAj/iK8MTb7P7hnTqtsSy1+F7V9zkyxTCZPBcjyDu5PI5AeRAb+DSmr
qMiyjv1A/Scxv92aUyEckoeLOh4ATUn2i8ipZb4jV0LcDtwOxy/2RB6qfUKlWXVckDYJqp/clAnR
shOQLHa8LDDaD6QEMEnR7IqX2HKohRDf/WWNc+yOguAVrmDHLRGJZ3quaSdQ9z5x/iPvcYQ83b2W
koYIug0dOkaYCtv06OwPvBZgKiQiaSEhs0SjR2JvACVgNeJLPYyFdMgDbwZ4sFo6teZ6IVXrebGv
I3oM6EBv3FFG8QrYAAa2EvR4HVsZZ5HnQvA9u8uZXMWWSi5EFUUnOzJAzjobsUqwyUEFqXqjy24h
kBWrW25SD8qfEv0FLqZBof0t+vAlxCN8wXHeJ7uCwFmJ39eeonO+8u3Z9KUlkebsFkJixsctx1YP
cJP1owo61eOc14tcSi5dCbjiItWbbrn4DzlJjRZuwZfVUBzIgtuhyAGXcQTmlOfJLdB3anf70IdX
GTgRAYVknNbyvDkYZooLdZZBrCMAleAg3zc6LWNb2xT5l1fMrS+vLT8ZROzdLiXL0ftgiVb5dzSy
mk5I1hfrolrf/bUR+lj5bfrsCPgkGgXEMaZRUkC+Kv+hFC/6w+Lwg/OlIf3QspR+XhQD1ZcOer0u
lN58Q6/KdacvRlcw7hOOu6MJE6njPhJdIiM9/BIDBRlemsBnQLkD/p4zRNunA1Td+PaxkllIg8Hw
Zv4hWuulh90jtf5q2t1ykaDipy0t2ehDfAbwmx87duA5HKODtZ+ijaXgPLzWYRKb2bsG6ZivXFh0
zUnareA2AysaFS4VPh+6euh8Nf/m8/y/+LVBCuZmqFv6wE5hBBo++KXTBAUHsKcTnJkhH83VM2OL
OjsN5n0DNO97ZDIw49uSHi2996Ta/3Xbd3vNMMGjPBvh6sALninxrhgMjazv8C8gzo5EW6v1o151
RHkjVGgHh1AD4t/yVWD7xtuxn8iR0KVyh5UxxpuxjkjsN7R+V312NiLTR/frEr53683TDlzNgwfr
2olowsB7BoF/aHV7GGKaaxdDDPLxoB+QK2wOYQUrc5WXLe5XO+mx0jI8xYIMvXN+I9rWEQOyti/P
45RPULZMo7n4hGA+opWgFl4JbdmeWulKWVXIdLCaOkOc3ty4wNlRUuuAn9FVttEoHU2ylECzg9fY
tJlmyAy7s8RmIZap2ABkjRBrejhX3IOdbBt4oluczMD54c9CWmnjkw3ebIS/XGG8mNz9at++M782
3f29f7E8F17y4D8X/wo7mTLhu1FBNMy514Qcz/RFJPkGru8HToePFmDE7AVJ2oZmEnsLdj/bmY7k
s6jNJu4TNCmcco4iKGwEV1pJJ+bXMOz48BZMVbb1UOSuHDzpZRbh7DfXhZF1sfR8tZOT+XX3DQZG
o0t/TES+LlkpVx288OP550BGC7MxjNL+jwuhtRaL1MTPpRLAAl6H6d9PbWAZ1H81a+GtZ1NYqsQH
npZLB7Onvom8NI2dl7ZjXpNndfkWlbRC9QhD5mJJb3IskmzJ3aUY9qqkyrYyFLNtIv4WSJAVNZf9
FUswgIiDi0nEkI5RRdOtN4kZYA5R0qnDRfvt01yC+M6KFL3q4FGEu1dwWEf1E2e+KvQ8TXtHOhzz
YiX1yFTjTjjWXr8L/V5oejSHRYBA2nBdxJrlAL1ApXAfsxmxcLF458EYTJewbTclF+A7HQG0EbXT
T4xb+ANfBZUSdJ2eLjwcAbijKZOrKfBaOsSA7QqTbdxvtFS8npWy1kMdogiBgb06F2RgNv/B1NAq
/q8VrFCEWz67MvDxPKz8SGnGYmdkDSRX+vTw9ZVAqRQH2xSVuTl1uq2ArZ4PI1kwKASUUBbqEiSy
k8wbjTEyFWCY16onpTIo2Qi5u/hGY2NrB0soVt+bPU2eTFKGPAXKnLB+p1TN++6c/iQkfT7+kiPE
6iAVwXiXKOPc+2fr6JUQHu2U68be/aprbxv0ie3cVKqGZZ/Biarc3fAZYcGTWl925vpIdB7uMyWp
uicjwWce/7XKKr9AuAczwv0tfsSwwhKIOca7g6BcloanvXxAuPRbRHJSHyhwFXfHTZjXmwm+uyru
zVkb1ORwGxchjMN0C1w4EROPpw8ERhDT7gxwrvyp5bVqtsDjYIOWdJQwmAWi2DnkaYB/p1EBdYiF
qzfzhFdgT9b+HNc8EwC18KH2AWOGRfIWquOyY5b7kIOImPrPsSTjrN/3Bq29mmk48DAx3yAj2bPV
9s5tQvn845tMPpeMgV8cqu4bkXcxr7Vfmtn4RcLDcAhSw4o8uwq0xgMERzp5QCx6lXH/huQN3GZm
XQIGDs2zj958UPxuy9fNxBXgxmgb6O5ybVH5ECzAqUjQVmczGdNydoWp6wMl+tzQl/lzhulLoUpQ
dzrkKVD4Y6Ncroc7VID/Nuix1DM9hoBUVkHwiisVwT9q54hKOPITExs+WscP9LkKvT0jsaJt5gcE
g+3xT8GrOg4Wu+O37hwEsZ/v3Ub25GK74dlWDY4oVyQ6ycQx2CTExngTclSIQPleON/MD0Gs8P3A
labAZaSTG2gHvncSorn7Y1bXkFa7vZBLmNaAt0v3I9FXEmGVsO34USnVlGeECALn3+zd73ySlh9A
DQGn0vTKqaHPV6gpTo6pwElAOz+/SFKVgHtkj81QLLBd7WupSgPTCO9qQgxi6FeqmmivxPM3h1U9
ojagv16dZ5r74w3WeRVFdiC1lij9peqLVjrViD3+ta6qnIc/zHLxtJmAOqA+n13adZyvGVII0cLv
3KoYv9/smCSsV03KaMn8MeWczwXD0WnZIb2ZoXLXO/VyhhljKaTBbtBWrug0oEPNiWDpPPWNqF54
5MW+q0E3mSPivQiETGRjRmPnjfAYkWzMXJcVTb5IH9dO6dtV9XINOzjOrel74On5/w9TmS0ZPA1Y
yRghJb50rtY89LhHN4+yqjYg1kayYKlC1O7v6nCrTw/zzdSAim++s/09Oa6NHLPaWJO1PNzNew6k
ehMlhZP6X0U4zB1TTG4onDDlFmHZa5sPU4ZPgnG7sZ9LpRKQJ1cineREp6Tje4k8wDk9MuAkJaah
1p6hCovIUELAhatBpBKjSHHZvML+Oy8IE/hWCcIfu37maFv6ayIBoHyUFFuOCKZ+p13zrybejfyo
MuQeqFbjgLUEbac3QVlT4q39T+sLigWXIY6I6Q/ohHr11oXvFW38K3TipK3ajG6xDnpZ8aOkxKmK
HNSZlDO/JOTK9wDWolxMDhJ4CMW3/8BRQqhwH+NQ5Y3ShrOMqVRdqI6eBMwBAfH8MKqkfsOXAGVp
oi61vuFUwco3/uGAgFgdjCiIJAgWPhR89/XgolX0LeZJTIvTDBc/cFYcqewQrTsVkLYaGav/TQO1
ir5fuymHOhqid9Mg3Gg9ndBqkLbHNgastOp1zQhaf/IRT6IrdDmjh9ye1o4H9vUrTAcPX7fiOVpc
LMqpmbY6bG9ImFXMv3goAxV3t0E+1XBEYTMEqMtd8LuCi02YVWHuiL+ilVHY8qnx5uIHBZAToLsU
dkZyGJvPN/9s9dwVEFltqBS29Oh1uEmS6D6jyRHX5RW8VfSJiZuU7dy3rrxWoc18JhpX2UojkbTK
P/qId7K/xe1G1kA2MHVLbN9n98n6c4toK1bHwGYudzXVcIJjgDGQRjl5O1+uxJkfIlB3L76BmnwH
2i3EinOC/84Bv2VitFxXz/9CK4yS2h7M47Q6K5zYs6V3Q8Gh3OZL26fHJkd6Kq9c/8CShCJonLbt
x0FDZL8avy73EEt4Ss3QKHt/JYuzG/TbGMopzWxT8idEXX62SfLRba/e5T3TkDaSGMsmHu2e6+Wc
o7WS7NDrkjo5Vw1mU+yFAmsdjHwB5/iNJdyhox2OkXey9NuJoHKo09ezGctMyrtCcyts6DYKVd4A
VxtvXSEID1H55nLz7KzvhShQCFXYCK/U5rBII1iTM3e5c0AqdkHU7hdNucMWAuVyefJFoTq0IRW/
th4z8nHjRpJR8jKTTXfDWdcObGC5qXKEFanHwKYQJvJbOdqT6Ub3jszOx54a4JZtFmI5u6XqNDTQ
Ilbw84tepvbql3TD84K+EiH0jH1Sn1/6tFYwx0xNO33nsyKessaWKYjLcTsW/BstqhraYnfqL37a
EgqZ5zoKcxMMln82wNwscj+ifjdFCVTyE+F80Qa6CI8DBdW+lJuzyynOCx5ZOeXB/RT5a6LZcEIH
MBUgBarxiE/kOzA8kdC/rDLAdWX0SibiImE2GRtYsP5PIAvM/MPYFWCtXMk7L/1X6cX9fAO8LrI0
6cPtkVvjnrCLr1WAwlfO24qQtdgneCIACqNrXckVILGsP/e4rnGhFKsTEcm3QpYrbrD5t6TPstZT
UcnTm/I/QAbQmeH5bwcDvUJ5A/ttXgx63g5axgOPW0r2SJxHhzitDkfqsBwId8JarXWWXtDjhog4
Fy2si8cRp0f4RWXEUS6KbpeFl0irdzLqkze/inL26NygydJu6PbQcXugxpCcn6q5dbxUu2UmV9kN
G1KjWoeboPrs4EXVBN9uHZraaDIFUNrgY/2hEFmIKnsBBFFPCzHmisF5kWsRJCatQZJy9kfSvTw0
RS0sPNdJTfLU7rIkkeHhkWGGx3Vh8OYqIf7X4Af1ItLyMZuAIX7Nuq7a3kwyKsbKEwglT/8SP1Sd
97DzcZDL0ejLaRFkmKQuDmkbEuqkn93MCL9dhQVVv3lk8D6gycukbQ0OQP1QGCETWZs0tbJYqX9u
/jj3RqXjDVezSUcrSs+optxU5uTONsRiAtWpOdRLB5OisM/iOouZ6hPzu4ScUfBXRK6SqcJAfosG
XVmShgTtc1nzyOsTpiwu4sjA34YEZdDnS97yHhjx60rnBBDl6Pq+Egws/v7gMVnwUO5/tiC3sp/O
g6Jp/ohitTgeithrkV89tC2/I3JehUbL/2Ds+ogBrYCJTvQklMxQsrXsVyHbVdlZmEBuS0gTXsoi
Xps5KA+rHehgyjeB8sW7LBs8Jd4+PO6q3ZsYYa2dU8ndL54gASg5oKKuWgcHpJd1yKH58mT8Y651
2AWoCbN3YUESvVZ8n3DexBDJs0roEnxYlUj9fVuQmZDdO/eAqdVV1Cq1ZlWnD5nHBsHeImYg1X1q
wurW4jUEvJqHA4JwyK0WS+ZW7RQnqB68AVFixDAcxUPg/9CDppiQh5TCsnZM1v6mKKkatC9OhCvG
/npFqp7i0gtpsHuYcIbS9sVseJMYwXAP8FVnq6ncvBlNwNtHFNr1NysS6C5ndveaQ5fHTuGI9DXf
N3XNyqnRdJ9V+Ft+9I+a8aFL7HBJA5mDcgoXDN+qyHgCp/n/vGcCMe1ISpHWR/QSjNvjtgOJ4UMs
+BSR3TmEYDPesSRl5TgST9foWY5XTqXTLHTRPWTipA8ndVk/T25oyZDMc84QFBX2lAP3II7lDsQg
5ks4cEUtfZfhvh49cL+lV1QTksIff9d6/t1ezjoeeDmiv9VnE+FtOm7Mfa5lShKW1DfyWScb5eqB
XtSTb8qU9/o2kKoF86fPS7bCxcj80mRlb0d+tXfOks5bsPur3oJesq6FY5WIrQyuu34ToSpWIAVK
yZ/J+1j0UWRstyzf2emQDA2IkTh6ZXqwjXXgU8NmEDVrg5KzUyQBoSgLy7Nu27oBsF9mgBl6b4HZ
ZW9SV2YdYFAHEZ7Q7dVUkJgWsIroHcZukcePr9UhchGfkFPdkCBAyCIVCNLWMwhh1KS3DA5uf2na
UIskTgcnEfM6GYAI8Cll/tGBR/j8rKyd3MWw9LtEAmbg4tIBbVP+gfVpnZmRK9uOsmVVMCIRzTdt
YEpF/PrDov/Fe2a/6uDbGLiqlpqgK1bNgcimooAICVqLdbs/sITFlfFY8TR+y480xd1NpGaYosK5
sDDze0Wg8JL9S3RouSAMbDkkOKWiB3hr+Q8rIxtryB0w2o18dH90DEkAoGgdorzww1UCQQTkKjkS
FlKwAtvGTfSdGedRy/f4SzDanMl+l9/Agd3zou0GAfYzdQgMoqzkMf3e2MkLcVRIcBvDFAEeeQhi
Ld6nnUq/pJdL7d1SV6+JpwApnYIAldjtLai8Shz8hswLKEwB1Ez5azOSd0BoObXe2vChwpJxOXdJ
Fi0nxJCAqYRUAi7g5/RjqnYIUeKzYXC5MEy32C2gLRa4L41ro1qB9FtM2kBj+qR0RhNxzjzmgfkd
qicINZ4xor5kP8Vu0snNuv4zI/p/fFfsjZbXBZOhVyWOQlFmx1VrfPt4fT00ElTsBUwr4LfdLJN1
rlw9OSptlnrs1XNKmUKsXUZHC2ya/b6Ky8v8/+hO4sDv0zQg3+IjrhIopcY7vGnJfG6zbFrPiALe
5uklofSmDdHb1LYQAEX8l75TRK6VmoXUPDje1isXQ/19iT+nPpjjSRLyhmxoNla82iBy5vE/pKcu
r3U7KahXY4pLod8ntg4V0JaCy0dLEzdVVaoI0JQT3LpNJEHZu+E6jhhgi5djPut+ysh/Cy4yW0oI
/qT+DMvdSGJrIeG7rISUVgqUS8Fg7jM3GwmlGMc2K9dPOJxPXA8nClVmx/RRoDGrc+aKw4uojaDm
09iEXqIBk1DG05JYaAeMf+0wgCBeUKg8WZtHElZroqg/OuKHMYbrwAT8LHoL0FSVYtzYdhf+PyA5
BWunYRd7ifa0dWTDZ8gBRl52uEIQTqCNNjLcepHn3YUiO/+WuvBtGziI9UnHvaAPI3mSfNkgYytb
I+hAJoh68CQBx5GrIOm1Uyyzwku1oQZ1bifs+0vSBaNwENJyEf8W4pN8WnnMa5k83uZElpjQE5up
EOdVypjfDTpNDV6DcUhdhRU20fgaKJ/ssNESCLPT+YzAuaao9Yr+gxlE72fN3QqVj6VPjpbhcSCM
hg8D+pLqYdHbFaDk0qtLuzaAWXg2Vk3xVCNeNhEFyJwvQe6kY9vJ0y50Z5iWbaOhTuUsJ1m8nfoj
BBNw2qjvDmOHJmu0H5rKILVSQkxC7TCBT5JrujuDK0modKX+54+0ORed5kZ5DH24sTBqhzOcqlnM
kI1/T+xtefDwInnrQDjQLfb0X5+MAw/M8nB+AoEDa9+N4ISU2BzwneMhh24BLjr9xdjvRoFRRf7U
e7M1WuZOvH1YzjFszAUc08JYduVp4/t8bWlhKp1+Z4c5raOXWkySP/bCtdQK//fKB4vv5O1YVu55
rDyPlh2arGiMVeybOC06T8Poi4pf3armR3CzretykkDuGusYWj79W5XapCfUS5vCTOJaGBI87I4z
8R4+s7TFnvpfEm5ZvW03s5ugpSb5r/OQ7uj2nQ8O5U3SyzFnTMBof3U5XDnbTzDxlaDXkTKNLBY3
wfRb9DCynuvwKbV+H0DQP7ANVslSkPNgVcvK+BFqwjl9fjxngqpaZluLOiEuwfXlJW1OXNFGJQM8
0aikXs4hq+2oxnpyg4EHycm9lI/vwDjaWwzkF+3Qo4iK/U20gAs06oC6uhd7gy+rc4hbjvK6YGpH
XL1ewBCe/WBWDH610aJGGixqYTfoCJ94a2yjhrsiAFXh1oAVZWnCvkfsTo+30ufcOntWb0b9qCRv
S+ndDVBEVg7FC5R0nCbj9FoJQC4Vy8CU2Y+MJ1nFqQH7lKTUNbNzN7JCmVpPbbgRJpHingY2G0oF
gxL8QX9f6ALEDrYg21mPovs3UK/+WeO1sbZC5htGvWFdiRIkBehcDLt/JfiU7M83+tC9aVpyAUz3
e+yc7t4qPtgmIYtOQCq907RcYwEtOc4TdcKazx/ldTj6s7/jGkF1xJntIjOKchJ+jmjLoHXUn0KL
LAUd4tGrWPlZdrrtw23298j2kERji7UmayKJiIXPYFvUnej9myvgADeQIozQ27mVG9qtQoZNkgEu
KkrZj2MpWb6LpMmO+4tean9VWxNnkXX1NTqdwSmJwBPg7E/rYvTHGmQ1gXK9qKW0zvYehuk8Hk3i
xlYj47aExxx0o0dLgJco2MRSv7sLGqzH7px0MS/d5OvV+UtEUo0aIH0T9Pdd34wKB+/bKzDsYewO
Q9IKlblF6LGn8IjukAeOnlePxM+YYlTVwrsxoNljWUeGKlMwZEH5kV/gNzlCaJH9sxiqRgrVTcK9
tezPKnFpZ5aI3ZsS0BwPbobrIHb1fV62AgQSC+paePLiRXI6VILqUlOQxHXMYh/o3bS6YxUXbSpe
kl5C/Ld6bWtfnCv6fgNevucmbnn1VY18zzKR5m4wuRanScMA7cL9w/wvXSE1IG6z5oBPdnDykq/r
LD81XY711Kyuq2sKOZXGzExQzQtZakfCDKZexpmL0WoNN05EROs4K/GnMcOypCDXUkF2PrJsTjTB
bDkbvxIOQuknEhCyFVIYsrXM5+Rb/rcv6r3fB9LMrMdBJ8inMXtCSf5UhE4IMSeinr7LEQmXBPNl
BSZ7B1FckO8APmMwQgiAsbtMZ+79EBPbUIMRAJLc7c1pqfz92fccN+/2VEweOd6zpXFujKojRDWo
YHODGH8WWa3+Lm9ucItCB/H7EZ9wsaRBQQ+3YGgnTcW5asyL8CkQt21ijkz+VwyTwwE7YMxOEZDV
gGMp/upOFSMDoMqUTd1ZV5OpoGm+yKbu0VBdAQxUeF9losmaorkoEWrpk9JltjOb/N8F0PSQsFf0
Kz6/r+sxKmMKdzRNHKs+VVNyUFfesh6/cfaPLxU/3ntTWVWRhtlwKAVCpbIZ3rwVmCEJgiHLefFN
+f6QIfzHccArGCPnwDs9Jk3tsG05og2h8q6o61BfbNPXYxVtkpY4TACb2NWhVDpgjPB6AHDWvN4L
/MCmJjReZVjOZR9zJedoQK5DQ2ZZ8Pb+cpW8QK9kFwtITE8cgw41gF2uLTAcHzrlAD8m5lcsids3
BEp7T1s4RnH1U6qqJ+G9HoCmp3ZUr9P3d58n/X68GS20RikYqrzaO3u8+y6tgthrRSkDKIpYXfZ4
K6qM6wG6Zfn2UlDaUIVrgkH5nLOirhS+bCpMR94eJ1RIfGRnoDgHFiqbO2EdKFe+C7ZfjvYHAa/Y
OiN8m/lLPBpuGJu6jAyri+kcYf+wKSPX8yxkV9DYTnTFA7Z2VYPfLSrmtY/NLfON2nxqOFJUMCpq
2tqIs8jrPgyxgbH2vQr9EggGlPnBmc5cvv5kcZYzhOwAemIrgfLMFbJbfkmzAL6CLkCkIluiTwEH
KBnbVeWElgV30seiVMEtQH5Dq4CYCX04Or4YC7Ic53HTW8cdgMsj0G5yM9/GTO/R/tkm/BInojCJ
9jK6qShTEjtp411AW0NV6Ux2zxn03t1vYCBg5/2nsHmRhXWIH1XgiNuT2mt8e+e33BNaIRjny+dj
ofA9VO9SOWmTr9D8JAG0rSanHQ5GnAnFvWPoGTPWNDBxmQwhxed4LKhLVWlEOvov4P1lgXe1NDqn
HeHhcSk1pNzTKCTmOfdKHGUC0X9hxYAbgMxLJWmqXAf5RjS7LrC7tApTOpBcKfVllT1EXvhMTWB5
5HYRP9OKfE6iJXkHmLttvem4YxRs9DYW6XhGdTsHEdnsgboYKKBsJkXClHcvv6ZTBB6QUzfYYLh0
Cei9zJQnir21SC1fJqtR//P3GL3RJnIVq75NI1PMCbNasEHG3p9bVnNqAiOeBU1CdOL9MVzbMDg+
RsbIUf2xgA5wau4QoxzOVA6ZTWFPkXYBrHvh07hlSK2FQ4JZjn/iTTwni4ABD36l7uEUSTkG9jha
AKTZsAJdKuz1GbTmtYXLPB3Dq7YW0TvorGRu3JvqyHlk0pE0UgwOVIt+srjmWppNG20UoRDQmqK0
dk1rpHTtc27R6vTjdvv8LU+KzILDcMi1Vlq5t3CYbybzjQTrpgdnllRj35yVDDWjxcv8NF0ONxb4
PAPu8oQxLjee869guTAnB4NlzaU3l1L6knUde/TwUcdF2LpDevWEfC+HGTxpiClZUtxH0oOSvKRN
9FzTK+BM0m5RdgW8Dqq952isjvCSi0ohP3J3+dF4BxBNKOjeFaG1Tyl32/FZA25O/hqCW71enZvd
+1AGriidcuDsPAw2/ZO5YESHG+tmcq1ONVDQ1W+NjZvjY16qI6GnArhTKYRNmcJ49HjOcmF5BLsz
EfLgEvsqvqtxu9YMAUmK69jW63dDnZqqouIdJSXiUZhlLolQUzzV1aAPjNyCU0a8A//Ux1v6f8gR
A4NyyR7XDsEgpLMm60cjYpTLvgtUCdlhnuXj0xg1ppsKNE2apsN3B94RODXW/AA5Yu17T6+ldicj
Ffk8dzeVEv8NR0T24FSuHHYe8dy1az7inmfjxduv5li6Yj3N9MhOzRl7lLeg2h05BWQadWIXPR66
HWEnzTDjbDlsx+VbxAouwY0PR4PDdlhmqPnk8FcW/ArxtN7VeeKqMmKs+qIKuvZZrgRswQEu99Ew
Eu307WHXwPTWVG02tmWERR8Uqaei19e18CldFEYDrpjXxO34rtKKG7qSHz4Hule+PCIBZVMpDJsO
fCxtC20AJfoKaNME4CUasatiUK6iXNauTEFEfRzqbsIlRLAskEIitXgdwsWpgDdOlhi62ul/dIyV
WHxFMT4Yf/ko05V8C9p9R5bt07SO0Yhco0tabGHmLD4Wi6uW2xqPXgYgpsG/K1QDOSF9h1K1+C4Z
0psqPn235S+qVkHCWwfZtYQ87XluV6Lxa3AsR6Ojf9h3SJfKtpC5hkdr/9mixyIivXE4/Rv1oUwO
lkk4dodT5tiQI3+MVnAgrFEhEMdm0kY0R0rFIeXh3amgvCnVXVTpmXezQKwwaByUP1YWv6/UJhK8
LxFYcSFFtxvIH5wCAlRW9c4o7Q2kyuec9QdflxI1eM3CvMXoXEW1p7MzT5qtpfJHEyeTqxwabubY
E8eUjAN8zdD5FUzYC+ESm7zG6EPqRfBW8DA3hEVWCIxzDjkh/vLMSw98e2ePQTlVVFuPQO1hcvNh
GttpI8SGtKlqDUHojTBwBVCO8Fa3+lrCOBZoYYkHFXxGatC2RRzBVvMH0CwQbhZEkz+MhIjDib+U
BvV/IFiR88qgIvJL+HZIJ/QmFHoiUo3sVkMceuycum0UKjFFtJlDGZ/DAAhLCRumjgPBiI4N2Dka
CfILSqQOaxAIKYpvFEbyWxGpaGcu9+06Dtym041mb6PaHF+jv3Viw2s39sJu9Hs86SuDL8qde3CW
YA3drupGMXzXW9lor8CgG5b4cLFtUa+rEwl5wma3Nv5oRZ0trwmobr4pGTcLj/udlhRVviE9/zP/
OL0j1EHPqqVTTm3uC3Bzie3DXyIrT/+f5cZ+oEX4KeyLBZZwxjvgnPOvgDHy/FfMDY3/4XLQCZUt
QIsZXVM6c/xzl8ujYW860NwXYsEeolOtyldvnwMhxFt6HL55NbSlXvpnC8vGhcDN3yNQzVxXMfQ1
0UpPzahegJi6iNji3mnrXHDC1ADTrILcv8bpu3Bd4YYr1KSc06ceqgAdBuxcD3Wfr5oCMeq8CDyt
9zcbmcXEJKipxLR+WYWawgt8ynD8wOz9l+WDDLkUxRB3Qtdt6VBweiqlOxo2CDY6sDZtzLdMJI7q
p1WEKuBMEhVZnd8egb+TtXQe4kn6azEqiWUTt8JLAd/mvS6g0pmCDxrSfHUt5XXGHuNzldsjxZQL
v+2SKkhKMV/V1vRJnnKkO3HhZuggHUDjTGRYXpjvd7kZho3D5IjZNCwPOW2Ir3DvyuFYJAq77FbV
87JGxDMjwUMfRecbXtZcKMNPKEHyLuuh7Qcsxnjojll/ja0lfKdmzLMDaCT1C536PlFTPET/diNb
XGTsrp/xutlNDEtqpfd5omiajJzau8ETmrEjaT5YKfs4f4dhppYAK/3vVPdjh6xgqydIC1UGD8Dz
utPw632HvSHLuP+tqT/LvQRArxN0j+9rq8HrWHnKN3YhFTvyx/K/LHCM8ZQ6kqjlk837n9WDFIQ9
du0cIi1XUk1VqBgvRDJxE2hb4PgwKZUh/aQMLPIWDZjpVVTkOBgKShE9RrYeE7TUwWPoOVUtKwrW
PcSsqIQjkAzTU1h8pPa4Vw+3Jwy6ji/7+m0PK1kX22aXm+HYzHkvkxWWe3JAGZgddbz3oeS9B6G+
1rZxP7YwknGgu8uz9oz9VzD5gqB6qJLXUHJjl9PX4QBIUEwCWFc0fiRiFnIU3AbZ9ZElBt/MF3x3
0/IuaRYmOodkTcW8UZF6FUwxWLdsbNJIEBbH2o8j4iOTjLW3H1sD8hCK4gdBEWMPZWathfcz7HPx
406V3wUbGKfSWWx9CEml6apRKJVPEc0TQp38nqSzLNIGQ5r5Dei8RJIeopVydQvTDZdLdEK5a1XN
1Jxh2RLkXQtTp2lb/YPbVJPRYptnqq6wqoGj9UquwQZNDtsugM0vFZVpSRErz8khkLzizESge1bR
U9NhFy1P2U561X2syaOI7mzWwIkWK5hXl+ObM1qM7Wn87xym9Xa3ELVWDPkeB518WtcL9Zo4a6+J
MpdytlVAbemGCq63hfiP8OUpv4LNFDkEsD529W2Z43UQCGmE7pOJSrZekxOuFAdwTebiAcyCpR3I
uP0IgJcgFJhNrtqSRp0hr5u0KuSx84v+zpbu7lEO5jaqLkg1xOOOiJYhUwlxeXD1/TtDUFxN/UGB
kUlICJvOJ3wVAaT/cOW0VBet6+7oElEW6982krZ1Qdtb5B8AKD6GUtDmP4KUM7rKp/Vq4JubYSbx
lalptHXv/Zw7zAT3ZZFwbsjmFUNmUf0eT1NmbqgvoqndkOrlxSPBOdkLXj3tfOmVvePvPvGkK6vS
yGoX9aykahdTFOgOOWvf/v9JFYuIDfe8r+mflgUGyq5Q/uEM+h/lJ8//BK5CxCY6mv2nn+hGpvZg
EbifEdO7mJqAd+kq8i10q5XshUPRZOxjghP3zjMOPWUCPB8aFHCyJ3REYVaLg7SOn1hD2DD4+aoH
9ruolVPWKcGEyT9eWFl94+22tiIMKBA3+PBUiCy6ggWeW/26/W0gBRyFAPFzn5ZPkgawX0xgtnfp
b9EY1ihvm+yT6XDwbnguiQ1vg8oLbNyN6E/JQ6ylMzjNstF+ljfK0t4ABqCQc5vSfD2ylXeWSrCy
s36/zIoaFDShJ57dpzG28MQITyhOQN9vM/3O9GLyJLRPRAjj2trzsJMB8Gi6J4XEZkFgMH2avKBJ
3EBHRTz8RqLOS87QJHn6pG+cLJiKHz5C4rgL8p1A1lK8YCeoQXC2uB3nDHx4+05i4yHoIGGnBdnO
n9VThMCKSoy5t91LFkCqlgetx47Mu97GPEpixE+J0lbl3siRyp++3Ub1zO9sN0CmCfh7zA33c1ya
ReMcPZ1dOUPRJt+U1JAFZoYoxIDrBKe35TGlq8xXKC2baxh5skXgm5pca8pDoSPwXllTk3GQtZO/
rEsT/zW2inmpplE7dkzqOR5GLwWqkEcCaQMO57EzQ9DaKyoXYGXyiLyaPivvCrEHTAH4ZIzRsVbR
61jZd8gxXL8argKUv9ggE65Tf80c0p9thIF6efF+sc8BG3ObieDFbfR+v45H77TINh5q3C1h0gto
F6UHL2IwTk3XZNFvWLbR1sv4klIYT6z0FHfKnwJo6pDPizqyEf1TQ8FbUD44GuygEXA0eO0rVyYl
QVAXglIqFtdZktej+6eeWgkpfTP1kPtyjRQPbZBUovLe1DjtnI4qJ+pLGndZNsudwynWzhLsrYiM
WtmNZKpFn06xakBwozSOAUjrUCHXmAxnPtv3pkVVTnWXxUum9fCknDrEuvtCzdqSd1MmlPMeV2CU
rjhmPIbptzpKTw3KVyHvDUoT32Pyz12tFyia4M54u/xffw3SZzL6y5lhYTCDpB5EKF/RApoSVjYk
IDJOCc+ayV6BRPXNU+LWmhSUEnH1gv+O0eWl/4ekTNP8lKNfpLJcC341bKf7lxE/qh/RHOCD1rZN
CN/UpYIkjf0PZ45Zzug86WYCxb1ExsLm3XTqNCxxeP/cE2lSdZJ0wZhOF31ewmypm4/7OQZox6Th
hoXmiGEOaCeJufRRM1WN80hcOjc7lOU+MYYOw942Ae4zttXvHHliycj2W9fusrSLR0UJoFdqeTlB
dCFKeNS2kyceLYwCv85dqjICXl0ZIwCq/mWTbOxKdY2QsQxGSaVvvOzyaG9vbE5K//I64By6hCwB
3TvzdLAmIBsOdkx3kCziczAWFxzV2iO6uWOL1mV+hBwqDOUM+H80G8Xpnsp1oaCbTJEkCpy9Luq5
tkHSnZh9FwdsEIupzX1LoE0krc7vB4lKZmkRXRVUKGnNt0zK1OPj0dwk4viiTiJ02trDEHAJED91
Z5ULjdvLxsv7fe8afFWD6qvkHE/4fkPfWdq5sRytYiYo0PLbw4suA5tKWSVw2ZEpVSA+q8wmyrGN
xo079lJ7t8bgPtNimPcK7NuiINkA45GjU8VDyoJS0XqTx1/9HyB2aOFRlcWO4eEoA3Gx3lu8IF4c
tl3i+iapwCLwSN8RS8zZndQPjyOr4Ztd0H0wJ383NegVViee3TxYprvblp4Kpz1FvugMDdZghVqu
31NJIRFqnagjd923wL9nvkC/Vy1/YwwU9typAaIu6uh0/kDZ5+KUVUgaFDcjJuG2fHrB5zfQ0D7D
wRzFjVVAWsIpDStaCjB61W9p2WYRFh7S7vIkML88OT5mDsqcfh1tdn+rikKF/c4D28Q0SluBDmOR
/GrT4T88s8373e8YfgPnJGLqim3CUvFXG25Vl0FeDlMCzUHjVGIj2wkyaI2mzyX2ITX5sQPaUKti
HmKZ81t9GO8OQ+KXsfjrlFseUZlab36cwFUMYxUjDg59ATXlAMUzVAEhGvnVGIlR54XXg4eJK4Eg
Z5a8di68wGHGc4+0d3Ll2cNxfDc1S0Jcw6neZuYjrncvEFhZqpli5KDkNWGO+1kXg2XPdnfkCvg1
Pv4T+8ObxWQOKFTGb0VOlikbn0ui/8wbLeP0cOS9lHIlzMH15BYsBx7LY07YiN+5thHzySZri9n8
XfymNrIBpIdsNH8xrSRrigiZurX7j/HE0bV3Qjop+o6hsIFjAGyerTWXu1fD5+4SFvEs6eeCCvCU
SOli1aRxIfqfFuShTvotjvs3vdeqd+mcFoCDx//hIQ3as1Oyv8KROZSEyt2SP5xH6GVTBDy1QS3F
fGkhd0euDRk1C8Rb28PO6pyRPmxI+duEJh8EhoZPmFRW29gnGP9I8vlhi79uaOZVU1BO57O/JmbC
5ghPoYkISclffXJqFbiiNdZF6OnVdnMQsZh7lH0JZJzciyyQeeKr9Sy/dQSAX0UBoK7WSXik6+Ba
Da1GHtqQ1uBPHXaSlsUCekR1GNAo20E0y+ZcdGx6Su+ShztX/40+M1XH461bEq+j9FVkuQ1a8X9+
lky2Vh2X7rqYqHbIje1kojyBiUV8KfhSlGgO6Lad85gMcZpeU8sCaSF6ruflPLsqLSFE1pPilKqr
2Gor1/Un5kPYlK3ZcDaSASA1fkFGsWl52n5xo0M/8icThYV7ZKjwE2oF33dY4/ZKt/Z7bg4tDkwn
jyYHIzhwZm5yO+ItLbs6t3i0o/D/tG99fIh8X1JQpbw9hjkVTP5Z22xP4b3ZrfuzsT78BeKdw6fJ
a8QvgzHsZDvdAHdOHH4utPz3E/r16PcOvuR0JJFIboMg5dtpocrk89O5Zh0ZZRs///MDg42KUvIk
WJxvxex1R7Fr8jlIni8BkMtkl8S7Hwubmxp3XIC11Ssz0/Xt8nXD2yBdb/alkquCxvnBy7jM1bYX
MNeuhCbEOq46g33qN+x5RH4E0f/59JtaQnVw0qaZeCZuo3G11PoeQt0oeTtF35rnzgJeulEEwojQ
HHECNelHbmKfR+b1KY7zlL8vZk/yhrJ3xtzk8dsHxqsWBjhKexswDZBXnw2u63LnzW4sD9nZ8Eij
eKGomcmxl+ZaQuk7mkS1m9woNUbsPEDcS16irY8keWuezLeIhsn3VNX8ip2iKzW6v+BPjs9wTado
llKG8lzSH24RGSXG3vCfhom7xJwlKr5itBjWWYDaHpsq8FO+QSp5x1jKSjQO969X/YygM/0jZF4G
2KUTNVlcqH9Rsl9H3SV8Au5rCBab6NX/terl7RAVRfSWdPfGTfWzhq+bM2X75wa0aFR8GRK4hBao
5ERyNAjk1WPkLVT3z78+4HUf0auKWXhFXMreQhRrry082VgFgoNN2bn9UNLFLgZSLSGD5kWYYqQk
cu/id+rGiEJ4BmPK4Z667teTMhvkHBVzud2i/ggmtDbLhcpKamA4qWQaIsLnZZ6CzoNIvMSSvUrH
7+fCK7qG2Lu0ZpQJT8SyeJ8bN/mCRiJnOH7N2i5kMwhSPuB06eb2oa5oTlEQ3cQ7gZhCk3EKMr5u
EOsL1PZuIKdiXLHNPE+DCs6TXlz5x4I77OfPfi8qOZgDLtVlTCqdxFCiKZEjqmz+nUW6gQZuhBsI
7ET/X9LZZX2cEIA+ibMC81/+zHz/d/fKA1P9ze3/QyX4LdSQN1Im7ZiF2XKyzGii2Fy+AQWI65+c
2RrC/jykTwbtJIXWw7bRAADdh0ZAgFVqJ5rMoYtHRo3VYfsjnjzCL6turpiCWKohB9tss8ufUqEN
krp60lqnTfOWiJAUv/9ws22bKEeypp2zKDsK2GMbfypVuXxeSL6jHr6MtDygbi49W3+B4UQrY6kc
VI89LPPM9PVkjTY/QY7p/8l/+CHm087pufPo5j2VsH61jbiRHJtOQ7XkmkNIfJI356uJcw/wBjos
6jPMSDNdHKBP7BxQRoaMX/ngc2W33qMJspkcO1tYI0m3Yx7c+0o2tqdMFx8KT8pBGj5DzhcTJQaR
kYrkngQpBFyTxu1FJ0Z8IcwCjwHb+z/yf7Lwzm92ardgH0/Sz3OVs3SQTVXeqeCquOBn8sK6D9Vk
JJtSdBK/jDatDR9oEr2cOioeDtupKSWlCxt0R9xFikpPkO7LNPN5rkNqjG7TavUZZwjU4c/1tvq1
EO3Ywvim65GcqeD0RJ7ueD1cLi+DqhmC1s4Cjbx+3u0UhnnNP7k266Q2bTH2USwlo4BKvlpR+mXI
/NN+XnuOU0buHgQoVUlmfnRCakDtNf90FP9EAxVa1cCCFmTkw1l4zIOJwIzViuOXtiLVyI+NZRdn
JMeTenQiMBke8exPoQWUUjoHOJEGxGQycRj1YpYZttmRiwZQwJ4Az5z7qv58GH91MZmzk1WIlvRJ
4yPbe9o5o4RDdYX3ncnwbZoiRqMPxhl8lrzH3NBE4PDU7kKk6IvL3R1P8rDyHgMjGSaAnpcVe+ci
dkow51duY/Ol3TqZab5+qLq9bA47kphzGLoZzXEGxqUNHdm5+EHvf2O4zs7y4fA8rtsf9KlFB9CC
QNts7vISo9TUKwDUuCkiOqTo1wxpQtkGZphri5HCpyeL9mU7EzGTss52gjBozMuRbhu0Q5tVGngv
TULHv5tx5yuG1lfxhsunoefAfF1rRlVAtTIlpQ+VX4YJJe4pRwlv3NSNwIT/aC2ViH90MdeqiYWM
UItB67wFWbATuskKPC7exroPyRwWEEjL9xIiUwGXu0HYUs6NCqqRy8H+DXk/nBTKW25/s5vUTBzM
ekvM9LadEVnbzlYb4vlfR8Kqsc0Uzs+y6qIL1mv1H0KfkBSxFBFcIoUaLNBqISib0HKLgtD4/ye6
BuZl1yOIizfgqrxGt54Kc3lyG+hInfv5JYS7A2IohicQ5w8BcKf65ULgsVpkPEqqGmlCW8C5qmP8
8QQDPFACxQAA821RntEAMELApBPCfKYo5JesuXhcKfEHCUiGSBor2XhyXpB0GlheJcQG4uSkokGJ
+basQpPhYnPaPb8i7l5eULfKMV33l6uCvRNtf8vt8xZmrDN0zpzR6gekCuB5JhDkFQGB9YFMxCSf
+c94n8/gA2QBasWoWXbSpW/yf8BpnU1s/AGraRNRoTqBqowYSFTrKYFSGHTjtewJoi2OSrKZOMHV
gjqsDbTv+lYEo4AaL4yjbgXDGW/uNx44uDoHHhXqCl8NnS/Hsc9Y9RPaCRPt/w1saiJIvvJf43AA
QF31aKgQQb6ZtzP3gPyymeqSyjQDiwa1unL9p3AiiW8/JsjicczdR3ZOkK8po4ZksgXyDCeys38m
SecR20p1xvKP8eQHDHCxO3fvbcz21pAf4/7USTqugvwolyRR1s+vll8Q5cx9O9VjkRkSSCJ+o8IY
wSpTHuBFZFjA4un8OCq0WhWkIJonmhZ7tysfZxXtuDEETmg2ybPBC4PFY0dUFuZLp4bR2XjVF10F
eljYQP0FrJXkpwA0V/hEZuqCe/pV43nyeYi8PWJgHZQGCVyG+P9jdFzMI36t49Kyv6ED6ridIy57
DJ/H/MgmLT0pgFZ7KYaLVBrMmElc/n5UGVZAnea915nrfoh6Ckd6QOAUIeKtFxl796ADMhZ2+vuY
4I6BzEYgKwkGl5cI8WphKJ9tsKavlPOJS6JUdzGYHF+RsVeisUw9UUNVjXRDO02VrAN9fMUkvkIf
8kWfPaL3x+raHlW/sV25Zv0eZzg4vRpRWesd8Hk5/591EZTA2frvWt+Ymc/YzA4fNHJXvecLzGO2
NcrDzbxHtW/7bQJEtHqWWmVR8+REPjZIsbFZNXd5zjFD8BcnwfocS5eyyupOJWSslvvkUZMJ61n0
BhRXN+cEc4fy2ZFEQ4a9kLnXWEcG0Mj4VAEF0TVKQ6vUrdOXZic64/9JtjtV7koNVNryNrNDSCyy
bu5BjCOwvFO/mS/zbRLVxn1rGisv8MmOhoH5QKWfuEELQ4prXuvawGRmn/cMfHVSZjVC9mpQLUzb
BWQ/8XoMyX9c+PP7WEihWFiU0DIzeBkwXn3ahfFs3VGDDwPQSm4KYRA3R0wTCoKpKihmljQ05Q8v
o8IVeX5J0qIsNriC1MrXws0w3pSDAkbd+EBFZstEoS17GR0HR2TQBjBauCr2u99VQ717BeywhWea
P51AU7Nxxj5XGpMiIeHL7gEjD/JWmbIL7Ppb/R+up0tBpCMYKXvYO2Eov8kpoX8KMquD2m30D/ad
LhiaI0Z/2n/9A3Olp3u/2+Wv7tYJ21CaQ8mDTZeKCwBu1QFHnQZhYokqVRDJmEOPuAFFPaz9NJzB
+6M6ragxyhtxr/E9PBKIhEn7w0Sj7vWKZCi3aE60XVyzk7zWOauvNKCFLhmBw4ofLIya8pNjrKMm
q4jKTz0SE+oG9FtEeS0GihqwcIBtxQhebLaIzQHCQr/IHmXfjSXs6O4jyqua+XZf9j7xNxsFzkeY
nVMX3075erNDW2mhX4nWC3mRr9QryDRNOY4qxX8e6b3KINrQSYXL/RSmB21FoznLZiuHkXGa/k/v
bxbVwPxxWKOQrKiBCnXkmmCFSpRn5TmE69YiW5U/jY8Hta0hGBwalzdQzSt4UON0HEWhVrWwxDVB
zn8C4ShTWdVp3bzinoIecJWmonpHkFyn3YQ0icpLfOkQmAN7XNKaPjTlBmutGMNjz0Mg2r3Twyq6
7LDTA60aEA0vLHwNY/nU+bbkNofhDRaGsCcBwqesmvHvEyrS3FpvkObhM2Tr7AyUUybV7Wy77+gH
G7J5WkADodr9WTQ4Fv70VBNVkLeWfBrVoOb6SRA6WKzWAgMkjBiEPU6h0nGQbSwMcL+gGWFO+C9S
w7BMeFfow1Tr2BiksK2J8PuVlgPO0wYdX+JLkZW6IDb1t0w2JXoU5bNzGZPTSJ/0qsE9owcbmj7R
hGnKZ84RHLnhC3dUTfZqu3lR4mdzi+KXIMh+3cQ11hLCd9KdgelBpO4QaoL1B1EQyWLsPBTT0ORo
JtRFKSJ+wyyl+3lnsbLVQn28Hn5F7mfNRzAnA4xhpsNKy4KbM3WcuptF0CVaVs/Jg/O/I8kqBWUN
fBHpYZBK0UziEEkvZeFoV+fjSPBUgvs6tpG7U3hUe2U0ykQhuIMpXAb5tPqflhKAuUVbkMwM3GC6
SxJx+IulFpQVlGmlxXuFelGbykhy4KMOKEN4nE/uRApXMbqIqxKq4jen2xsR/IXwLJhyMFXHJo6A
ArvePYbGaFQRtZ6OBa04IumYDJ1IkDs4ovfX5Jh7N2GRhZladt1NDeWC8OqGBEvZ3UIKqIe+sG8m
8fRmZa+JgVQxqaoADpjt/Ah5BETA6Ad+g12IsmxAPxSDgzLmlZblzwyozfXhRTL0+F07SiLLdeJa
sh8UdrSe1HaTwf7Ar3YYUdwJWN3hG+4DV/jVlAXpv3UeZ0ZVQA58S07Jk7l/FU/XJOWO0wjmYJ2i
y9V2JO93ghev5AZD2AxFvVn9GX66ydEQq5mz5Cz9a9CvPY7u1d7Zn2BHgWsZYQOp/8nvdP5iz9aZ
pJHFMV8zs8zUaXEwq6EfVMnDDnP2B++NeS++H9IvazY557XuWQ4+Lltt0/cUqzhgelFy4Cc7eh0w
c+mVD4daQGnShHrULcopO3vWauJQQB8E2dMRKGRcJeGwEF9EA28qWkU4jMjLxhnxzxfQ2IuhM0N+
Oau0CaXHzPrv8jTNKMKbC4NRXkZkWbER52y6pcgp9wDLxtdk6QV/qUoKFV4Earg2zo8q4/N3zT9B
hQ7c6sPtvBh0D2ywIVwtNspQ6Wu4GycaRTxjDE9/BIVn1W4XmCVtWk1IRhT70yAy1nKGOzm19QWf
qUmdAvkrJzr6Z1bvPvzB/Oq8GF7DwPjVfhi9GlvBdge7lCElvaKH3jdhRLOsOALAZdNHscbGNS+k
lpMgxxdMLSa7kfZkkJRmziHc+JHFMNxTJJjcI0aai9NbVUBywcCAYrHSvohP9qhx4++P6jMkRaoq
VwXU9JFL7D6mbouVhXmYtqEEqVOfQu5MMsyVBfHHFqJyIxgIs3xm5s/QmGsdhuCbgbkOFj/Ub0Z9
F9pGJKO3cTzM3zpzx+2djtCE0YdZE5GhY4XCj2PLkWs9Vf3plHf9ccwWI78gK44aVteYfXyzPGys
Uo4koycAP7Re3KwaUiBMQZSdA11Nv7ZCCg4C4Byc4I0obHDfXY2HvOu16fD35XQgUBmg7sasmPtG
BuzCS5e5dUXbil3DfZz9g+gHLMx6zyswge0Ket3ST2Ha1X6Kc+Q9ruH74LcN4pxNFbscEXqzfUNw
4xQkmZNHrLweLA71aXduuuPhq+34kIWjPLYVMnVC4UoYcq/fWx1EAjU52HOKI4M1zc+FkQX4iDR/
tsYSbXf3gf4By4tdawgfiim30YfvPBovEVzm8r6Y4KfQLQMqwZXbxhf3lvjHV6jZ4gbJjZOuAAEP
4LgcDFSSIaORolP6oIoGvWQ9zU6MGO4cS08Te8mPfa3iEvOLDeFUqPFse6E4AiFSUZVR414F42iD
bYhPxNkzAq+LG7hzsC+d5VFGp1OKtJNOF0HZPP0WBuy6CHMZjIct4kXaCjVWZv0sSWH7xb92FcpG
xZzTsT7J03Kau9rlFcw3ZRnla+sPdlbcrx9qU3bBNpaARH0w4cihenwRbEutplfdWN7UYrxcIrBn
0SbugOluUFbOe/Hc+c+DuXvHvWiT/AvIEjO/9GfL0XxWduLljQbBNQ68bw+rQBPc+E+pw6MHXone
4v9DZQRIUR1+6pLEwpYXuC4qxYGn29c9PU9074b0cumSAHyxcSpooFWd6EJWsKKetq/mx4bUFKNS
LcLxmBT1d2IgJUe0WavP8+nnN8dTeNah40nmPE2Hq/uQE/tMEb0LHOyufLYqiPW5jibf9KuwIKay
PnU1DxQLMf6p1LQ0SWs4S8szIEUIVdaQ6DR+wQPG8chsLvXPEekf0IsSqnvJz7sbx56Cvm8bIUb9
rSr0WrBc60HrJbGgzeDaZ8SSw8+KFl30KY358XwAhp46n6FYjC9lY/jbifbescQF1M/RNefyrRiq
2WrkmiCfNXqYfIlQt3optaTy4sgBlUzSsQoHPrAjY70feJjJe2O7AT0+BTQAeRbvcG+LTKmDRAcL
dP+CipObG21L8iF4kWj7u7Mxbq1WPC1HMj9AsisC2TX7KK9PJT32yJ/IKEWubm5cz5nZ4M7gU3GB
zH6lKWIGXnxgh/zpSBp+GVdp1U9k/njfjjOfO1/j4VSi9nrDHmR2kyHOArH9tcA5TM3PQxU68QdC
Dgs5wKMJzBD6xP3zFU33HxDioW0Xa0ehjnRTmfNd7OoJY9vlby6LREYhM2n8YNnauNM3UclTs6+2
4pItLIeKcyKxi/fBO7R8hPQOF+PG2Nj0d9Um89MwELpFT6cbwv6Uy/AUVfAHtllAwI8yQcz7roaG
6bWVCMYLnbCw5uBy9YbiArlN1Yih0mb4rVI4azaTeMnd7EbwdPU+q+ysYzilzX7IFJVGgNkFPzKi
SFoqW4UblGvkTc938bTUID5rDUjEAkx+aXMptbBxpIiP1p1B8ZJuOsi/NhuArfVlXCddtCrLIKLq
T8jB+jzkbB+24E87+Hfx4JzqY2z7T8sUq1C1vndEgWeBmLnHjGrw2lkRpwuMWXLmcxRuo5rmF6Au
QhOQ8nhbY7EXcKrL0khl6n30fZ3ZIXHav6VSVeEfBgWHHgAbdxcM0xUSIqfLp5CnnnSml085P1rl
bqkylf2LbcueG11Cm4sOO6h9JJF5Zqt1A3+W/9oeO/nvPWfHlLtkPsGgdHZLL/JIA/vpuPLG4nDQ
kTh3qzMOPMxkqHLWEvpOgxeUhBrTtvIZUL4CW0Jym5UsG2mlrOzMmbeGU6HBVkqKNhRtusbpL2pW
KccazJzbIthhwQtauUjiZVE01dCfgBUyvjr5Ze4Lv3Pd7kimDlkyhtKPeXsmegmKCOQDD4OY+wCX
m78ErofiX0b5ruB7rsAHF8kqIWMn5nJBbxEn2Vc/6utqcddQ87KGYcE7mtxqqzoxKPeD1wwPgv1X
kKhXHWb+Id3Gd6slHmbGUws9wOWCC1NAs3ppyzrJlM/QnH9SN9C5L6WZbxOE1aZbgTadQUJEYSzS
wOZA6qK3viYynvi5mQgtg5GMnjY7Xna20Ser8XEIpd5mp2BNa1Se6WYlkdAripQ/TZS7XXHpAKaq
WcEs2CsQxZ1N6Y2me6eubKSd2PRvsjvQCphxKiwrByl2mr9DrufcGnsmXXZ6uujDLxrkkSUIcnF1
fLdqdzQdpQBwl28U6AZokJk/vew+LO2x4NmltBsPMUOzqAZmDKreCTYmhcHwW5OzavGwe5HqU5VW
CTHIO1BQQ9LNRTrz9gyjGjuc4qfluFi9sRYXBStJNCrqYkY9Jm+5LfP8I9k+PaU+FLwMX719HJRi
MTkkzUjep1tx/ihB3dhB6gX8Gz1O0/X4xv5iZ55x/aNe2BoeMJyxY3G+w3i5/4yvVgnW9MHVd6O5
y2Dp1a4SqoVaglJFQfE86Lip2gq6BlUv/ZjtVbIEGfyfgYxb+DVw/iojviLJWYep6Ms/31b8As+B
345X/5v5C+aeDf4n9JnX7X5WqcQh3DGSptHuXiwTPbr9J1mb++W2+ZdzdNPMYmx3rzZ3/rrSbVR+
WL2LDcZjhahbNs7boupbzpx5NWEKaeWMLporagFevh6c+D24W3mb3IJ7cH/JS62ECrjkSvHLCKdR
Jvay/XJ9FyStHAj++G9wyy9fzpGbI9QD+8VKqt50fxvDVyYFcz8ICNe8UjnlcMnqWyqtktKsQRVA
TdveM4JCkVG1TjzstjwHWEIpNHrQOm1x1NCb+hzAD/Yyq/IVT3Qj4jo6A+ga15f4iQfrmvsEElTR
nS8DWhhzJFWmpfTZAL+qqS34dH6v7Ga8FIjrWOdraRvChroaTAZfOWKuJve0HUnMFH346Hz3+7A9
/8/I209OcZ+p3FovtfYvh3PTFpJxSc7rC6BxJ+7edKTwDnpmx+sBXJQ34OfNfOkjeBaTI26iAoUg
vmf1uuRYMnCddRl+phoSnZRsf/ApiDFYvllIBTFfKJ5l0lKRfa/9eJ/Hr2xgGxPPD76MPlTZrzsO
BSu9ePZU/GTD+9NXgWrs5XiedlEX52wOkWaB6gYPHheCW4Uef5sc7jE8IyS8s3r3A8gSBjVAWVOM
VE+M3ldqjBL9k4lYhLYoixz/Nv8oS79Rk0Trc+bR0h6UxuB1iJiVhABjAc8gJdVCFU+ZFAQu9ajw
IUFVJ5JOUssfrlukf2nHfHjkK/ksZg+642cYF/DpBXGfVHzdsajJHNnYnz9j//Wh/c262nXIZyCj
EszYTnGwOOESuVkeLfQKoMUnJLfqBl3eCR6vlCTey+cK/CZL1HCv9tFML1KeARMQsdVNPa9QHJ8w
+7/2Kq2iAnwRzgkRwwybWRbfqMfgS7dO1RCL6UqQR2LTkvPWojrE6SIaGs/WWf1x1jkNYSp2e1cC
/YsFPJ1AA27SLYhurQ+mFz1AinspWefdkYv2MQ5vyjL/78lL32b6BS1vKuAv9MQjXB74daW4qr3D
Ho8SUTV2Md2dZ0J0ICricc1nTg1l3Nrpe8y2mBn09e78/TYP3y7F1/nRN/eM3VuSEfXwYvTYXrFO
1BhPLA0KU4GGcn+noCTbtd/Q6nNVyYm5uNTKCOC4O2hPnldzgTGND9uHUSM7VVdpVt/Y+Klvsz8v
CcfIqZIZtC8hYf4GFVG9XMda9jb0Zk6VoEyDutluFFgexK4qTFYvVq51XXonINtFNiAELHBBi5we
YhzCcs01k1O5DUWoZK8rG/EOEoYpx638c5vn8vHPGJjgW3AWT4C1QneonspPZdccXVafDsr05lp/
UTYC7IaYAHk1BIKmMnuT5oRXL5Cy3/NfufLCvMFrU3FIRaEHVlTQllc5kHRVqbGDzH+se1Xp9YPb
gcIiSQIEW09RpGrnKtqFrqbrftk4s46s91nHAupfapZ58KGIcf0A/iUfOEdUNTmi5io1LCb5RFIR
r7lM2lU3BzWxvI6weRZS718wa2ZfACjSUxxARwpdnVKD/3QAsDC62lQKrKU1SlwtO29tnLYHPlHK
fzZJpZpa1cWY9aoV/go9D8BTkzZf+uRYFZWFr8IH12LU9DVXsYY6jpHFiujN6trYseY1Oc9SaVMB
CD2ln2hl5vuhsKwaIlf1ajtmFSSqqTmyPbdSAGwZwb0itgkVJD6CPkoZwKL63c+bpH4KHQzXeFDz
t6OsQWLNBitrLiCgaPcsSGD0AYyHWwCM2ElyUdRY07fsLruPMQsNlbdRYeFhweaXZgzQz1fY5bT2
QNY7JtKlBx4BFmttjvMCqhYl1xrStd3KsBmOsNL1wWbd6u1trSZtN6oMgtZs6yNbmirbTKvdV20k
ZAXaLxPqOTuHB1zYB8jMA6pGKB8+Dc46TDp71Qa++T+ilXlXA1TQuvsSYlv+eF++H5iS+DSckVQ/
DY7O0r1M+DmA9N9F8doOV9jfx5Rj9BOfjHTEHqikRQsax5s4IQjzipnYRu5S+T6RWUHYlS2fxhBd
5Oa/m97pUq86//v+ClQ/4IiH6J14nlFw4soSQ0nxha5xgvJcvrNzlXtSnHjkRwhNBYfEhRsl0k/3
h2pLEzweBvbJEfX+0G/VCOETo75xq0y8yjXGCKob2U+tbvLzLI2Fqw7wppjTzrotsOPLZ5/yRT5/
GYOwLtb3w+881GIoq62+xEuzTWGJjceHsada9KoS7/q+tAFLLlAcWNHFoqR883PyjAttmWIN3LOG
/SR3Lh9t+negOoJ5US4/X1BdmDQpSIx4M32hfpiKSYia6s25RmX/Te03+nPRr6iuSYxXTiwA0BU1
HXbJnvefZ/RP4+25ga1WvD7cc5QKhSCPOWyQCedpDdyOBUykLkb3i1cMFcQVWDSDPZdWKfZNqQGo
NIOqBA/iPxeLypm7yVO+77aaCWiNhpyoUJ9diWrGm/Smxb5JOSQaK6g5/GbVxJBJO2ZOGw48QdMf
43Mz3Rt9wbqHg9lS9sF3UTjMxJoqHH7iYyx+GZpoVkgLkCBWahQA4QCf9GfrjrgMhmlxtmba7vWz
Tm0QkFbFKKEq8tG0mikiqfCVJDIcO5QYBpLI4dDBzM/7wMdpLzwe3RDXA25c/7gOg2dyYLjPvjJg
O9D+AjZHt9QDFj6k7j+IN2rF8Av8NY84nf6ALHSjIst1e0+HFRGt/aN4T2QlQbVnd6ZqaWLnBsLK
On8AgNpMiM+8k+xdUacnNAhn3TXdrvIf3NSouHKR/jWlD37jJMBmpZjV1GWWL+9Fq0tQZCuudc7R
JT0RgFKNOP+0n7ICWxWK2Zf65mRrEgkwsdoED14RyZDVNRwzQQD93Xex+iFEIcW6tOhJgDbIlG4/
3MwvLZhwMSn+qhXXANv6UI5QfVojUe9RRjIzk8YQw8hiY/jrF7pnFKRDm3oHLfV7Mv8qVP0wqivW
ogCc2SzopaoLp27Yy1opBJtVeouJaUON1qQBaIvUL2NoDStAX/CKYfVVjjTRj/cZxg4oB+HBW6Ed
s+KN3ctH1Wl6effw6C8HGSvc925hWzbkcCYb8K4i0lFc39VF7EU9lDURmh5yaNBIOSdXQi0vogCi
EeJrEXsXV5JMwWXiPipLWlFdaHxbXcVOnoni+yF6Sb7E6VAIQSOZO1HU/kJMQVUGRySMFx+FmR78
m7+rVukTYuU0OcZPP1dkFWEGvFMegVitIg6VzcPT/ntu0EdEQA8aqO0bEXTSjGB0k6OY7p11SoqP
cd+60NWf3WOA0MsxmmHUNyBCubXUBK1gpfjSwF0ozobx6wRCFNKhi09NNA3lF4+LOQZiOwVwS+tD
SiNvfWPtWEK2Nc6FQdpVaCMwO5qRDGN6+WkNMCavbezGC5gy+ELGYc5YEa048oOmStNAds90MNjX
qNQt/Z6DPHtPD0ejCTd0PY/nPWtH1E/lQR/1GD7YJzWhZx/KzPQfNH7D/oZ2rp9N62sUaDSgTRxK
/ulir9nY3JV+jeUol4SWPZdeyxX9CvD3UD7B5u6XGH4rX6jA0kIQgkwVtUieRAZTiAYU4ZHoaL7W
BLgkG51ySLl5wwgTXJm2M+XhWvHnB7JXvUgmOEshcK3yW2od1FXllKEn/+ruq7DPAOaRFKORorkt
JeN0H1gBp6QU4l9urdp3m5WKWGqCp+lEyxQxCwzNweqZiv+XVXYm0eNRuIErYO3K0slJx7IlBIx3
wcK2EMaI0rtoAZZ99WGvNDN7xtcUrr4MKeezm+bn3c9cjONXGgDRgdTnnHR7qBWe/6UGJx9Q03yq
bjklwlNqGy/cofqhC95d4lZjGfI4IfaKKYFuSC2gTh8zCMwEdKm2IxmfdcYYALWIzJYGbNpVxyXN
8Bxwge/p0//WzrSO6tjf3YOcSzkNx3QrPDMZGos2zIduDY/1DzjaDT+NUFbUXfbop5Yv1mluzkW+
czPVydRrWFw5u5KYRwN5mJlE04vpSMiyUpXxpjwcB3ME1ExPcilIc0JTKL669NHIXKOQOs/pcy39
wn0iIAc8ZdXsycWTAQBxzf3BtYZrUh9/Gn9ZkHR79OUyHIEwNVGlenHONKBwYdeurLsz2alRQPoN
vKVfDR2CSmx5RAsXAxewSVEfcpdDPNilXc/gga0JsUH/tvj0mALOA456BAwNjweRvm9sOk4uqzs1
iapu1blILxG5M8PpXtzXn0J2zWT55R28YzE8EZ9ORmGn09Tyl4kxkfJ331jEWTmPILofkzAVN1GK
JACv7hnIhhBZG6OfwQTPkjvEl4IdBCa/MOVQ/V/384ssCfbyhwuzz134YhSI7KWTYqsRslnHtICQ
TB+E2lc3Nuf2uwOWAZDK91eNTfx91QgDyQc31UJedGBUys549M/YclGDnCTXFDhlUKLLt5+snLCQ
D+rc9iy6SOXV/pNEPdfcvAoOMyGyHFmQYP6svyMIEpPb/tCXZvV9Ifipy6jcH9+42FM5SNVS0ypX
uth9C/kS0Kjal9uia5eT5X3pWSy/SMkKTpEhEvVgxRUaX4d6BG/28IRBKie9J7wg3RX/fbHELItL
IuIv32PzGkhg95jcUvMPp9Ctvjr2D8bUaj/Mtqnb7kRfjNv9bPaNjDZgI4Ok4Ia/wnhCaAhbf6th
ny/wp2sTsY6f+UgKPmIhextXaq9/GPeMl44OfpDZHp4ELPHnxQqfve2irL3tyRKagFjMAMaLADWo
9R7xRHs9ecZLYfrOmPp8xojLZ/erwsO/+YQrXS30nU8p2+ouD0/leTzKv1xTv0/UT27qyluS4SG+
wiCWIL8wrDtN7PAflm8Hu4wh6i7wOAwGX8y6hp6/0X9uuIstGhgDNTkRjv4nINsnyCWm/a5B0f1Q
b1ezW6SISX4MoV+t4j8+1t2h3P6xTHoVVblNn//mvt3x1JK+yiaKve/cqjb7gBfILJT3i/nzTs7M
lMSHVk+yF3lVrmdkkbv69efV18vqnjiAAtxE4kkOGVObQ5TjqX5Dovr5thrqIp6S87JD1efJW0w+
3lf1S/KKrPNkIw+x5xP4ijFeoaIUGmZlBlLRIyj3JYzcWROayWXFd5xUMuiyFpmpMRM7t4UIxMNz
AuZVVcFeQxpSnRQ+uzp1E3rJiyBdPeO3kIgbnxh/e3KfjEdj40I14qDwBoS27u4KVzAXCjVE2lL7
ziYkdAqT4oYg6AJU/y+CDQD1DQBZWdQ8TKy+cxQALgKvkdfUo1CiYWOSCGhW0Zzr6R8KwLbnnlNB
CeyASaW1wCkKjuZvkYIHVozU8U8U0ZZcrDYf+QYMV82ucUZV86Frr37rd9wWHuopuC/JaH23gDCE
OJ0IjlraRhjvwOrf3WjWTVgECxvOQHjgtuzd/6Ye+gqaTBmae+MryiNMYkxEGiZ2mOjENKTGWXmb
BOp4I2swJwnqbhHvodumSn6vpklC9K2vWXz9zAwEi+uBK1orQ/3ZkR8e70n3DNPsa6BHQeZp7284
5+fXrfrpJFKKH0720EPgKiY8N1P2kN5X3/Yc4lexTWkNhc9Kd6sAQclhel5C1yY9hg5pnMwlGxVU
wMEcHCO+iBDSy0/4TcdXwuoy2C7lUh1FxInMvYm6/S6wg9EOrBeqVKhUlp12cqw5+SWVpXFwD2Mk
UBOSaRdj53iUkO/ssmZOfpDLczJpiLTtHvW71AUY/enSVPEEvkCSWgZff6K7F/jvSW0D5iEp1LmX
ahpW+Rfp4xlBYmYEN4LvZTb//GZGG6mYsGROjRlet2oChVWPc7Fm6Jn1UYgfTo/zBaHAkRWHVLHt
GIv3LcEvJL6QivJdk3b2KavPvPUF8ff7MSYPK9v0Y7zASBvl1PPAA7GNF6n2jZ+yuCjDifxKmjbY
vxjsq1AM0ReiltQVH7QOs/TNFQAMnvV8uiYHeBEmrVmQPPdBTbKetroCbbYZWhLgbQ6Uiq1bIPPr
l2v2jWem2QUDZLVj6dlm7NmwIe2Paga32NeKb8zBfx7mjVMrhekHL/c7Sf7U238sfIgRQjOFYVLy
VgEYNTe5E95vXSSk7TDclsZ98izRfwVvK4pJdp4ik/UNB35faHgs4Zk9SqR7UIoOhqOhqpnCvtID
04e+ZSvlu87oU/R8JvqEi6+AIMvHWuUlabZY1Tt5maXKdMoWhIv8XHq3RTAExz8Jf++s/504oF1y
h1FUiyO2Jdjj5QTc1Sk10A1wtBc5knNI3IsSJbpH14uVtb7o9az39RPJd2N62xMhXqcuL/aNVPnP
FZYNRLp3MMgEhJUoCEvSH3VWiOgUVw2DvpR9AypjpVmfxVDDNtb0msPuXZyRKUWlnE7m1k1sXQXT
g3/qAMhs5f4lyySAww8sXNZomKIn1hTpbpn0RrF1T6+TCSyEDusBfAku/bett2AnOyVJW1stup4e
rYKf4jwM4XZTrU0mLgJQYjPXMcBCtG93R8854ncnL8q9DZIAtpZvbYpX6iU47Do8EpNFVEEN1h4g
02EXcd/43A7rTNjL3HZv9X7eQt2keaBkMeQ22BKCWCcQmgGzqW+FjUxn1ew/35GAHX+apzlFckWe
g9ZVkABnehEoCU8CLzmmtQHwQnvwgPFtO/C4jF4+8479rAv52+d6KwG33B0UfM4jwKmZvYpV9C+w
Ui3DL7PYQvnIp4dW+r0Wt5HzrHuYUX8z8OaxRMk8P8WUSmm9dW5nNeoU/soYPhH0VOINdF+P2fOn
MYURmpSi5PpHKbPm9uQBC+1rB3kMd4KS3pTmIbsxhXgSeNRRQpVyHshYnc3x9K7yCuku3yJocMfT
GsPTcGJ1Y9vM0XnjIZjkZT/SunTkViNPTwGl2JKP7XhtAexyTz2q0d/iGSyDh0sx7UNXwT4OSuHZ
31Nq1Ake3dUxAXtHdBdmqbA9v6P3aiSm9EcZj2tNuCeAg6zIb0KFq+ZiDK4U+aBnsiI10B7azpYE
f5OQOVlaXtTDVF0RUOCwDBCFAHT9rQYp/FaAOZd1yTg/DhEh/2e1IgmWAOhw4iOQ8uL6swGPMDMk
Qk6FnfynDO7qnQPYRsWQRmbmukDPVyi3WGqZzynFAZCMrHo96j0c/9Wgbs2gMVm5lHA7lpFaMsPh
FTGbRXb5Sqf0O0kkoGLQrkretN/AVUiOFb1Mr9A1714fqV4khVVy/l4zIqYOlF9axlPcTv1x7f0Y
2RD+hwrKD+AqDjVWyouVlLySjvHX8Ifm4Z1WEwUvxZQIa3aSDYKQTTZEKZwyg6nvzd+rG/R7YJTI
3EgSWucCkawxhDF7UKGXt1ziXmSd/WetSBWEdaxWka1L/gycqjm8hfb9mWLLSeenmdcegCAzKRfu
tXLsnaXVDoZ9PuvbEd/qp0+Dqg6pSnOSMzcB94t4THcz7PXd4WAvVqz2VjfiWWeGnzZ6wym1ySVa
MYsFxEx6qPVWRvjcWmmLUypgM7bHzXtMhnbHj2/h+RZg5cSgVay0enppxmVne8AXK1wwZMtuS6kd
0lX6sUv6QKnTMoLpb/vTg1STHBA8/P8BN3o3WknJUnluFkme0M0CXoiytnVCTC23p9WdpLQhOmhg
gYWZvhdviFcYmFgzbrFjcDIGR7+iL9n1vaB7TW8EeALbpmNOrh0psv2qr+nwMSQuB1mWy5RS/A3m
l5VQ23HuzXxZkoIC5PR9qpQTFf4PnRrwQpuHQwBXXU+2GsKwIacx+vsw+tydqBWdW+pOPxnsE28x
QJGq4qHgem9RPVHKgIXfUMwxtQSjvdFvxijdD8ZU04RGuXViCNT7H2a2VJHaixlk0bKmJATkSVn8
HnjoqCaWXe+x/RrJ6Qh8zZ3GFutpZ6lNJqsVsgC3N9H8ZpQzbw1c+IU5Alh++pqn7RhDsZTfzbDl
3P5D9rDbZU+Ar2wblFKzx5FJimdJW6WzEUtdenNZJCuM3G7D+FuArQuADi77vr/bo9DU45lNKIb3
NJ/Lug9m8kC0awcxlO7oyTxd+eg+viajo2QSGuTW7Ey73daa5MdN1ToST3Ch8Tu4R2qquRH3X42Z
NFguCn1/ICK6VJ/ol7DGAtIcBbbd2aBC+uzmlcSaUaZMja8u+otN7jciLmmAGKLGzf1/NZpbL3mX
nrU0CsVfeqG+WmTp2nsZzA3LekoD8jq9oONAUoK4xN5Kiqf9FIApPR01FvL9PSZojITdW26Ccmuk
Ssr2rwmItmln/+UqVtFDdD7hIHF9UkM8rRzdb7mV41tt3EE/2dc252i49FhZGtG/yQ3ZM5X0qASh
BKk4WK+hlgh4icAajYQVco8lmCoBGLf/4KhnAkEFbjkUecXDmfZ/nWIl2FG0JWhVPTcmswZ4elLR
2iLtN3PaWPf2FUcQrtsLHZwJAM5FBoUyFkF8LBAD9+VEnYh5gMP5UVSUjHcpgAQnkOsvvoMsfAw8
xlJ5tg8bPPCHdIzTO7MnErLr2vcKpVQ977fCD/FFVF9v0I+0zHODXk8H+G3d4K6Y0vaPF1E4JyHQ
ZdlXk1+vfwbYGUD5WZtnuJBRHec32zSb5a3MZz2NVHUp/052dmrzILzTKYeswQSsh19sppMgnvLy
jTKVE8aGsvZzugNusGGJdOtyosCkljMtpfIzQPEgGAIOgvDIOGjNbuzDkZRGqHiuariGNMRNprG7
PQICv06NOzPDK7iU/kKdzSA3OyNvUomG/XZpaF/H9h5Qh1wGwA8S9iyvXYdE9kRskQAVi4gn+UzW
Fiy79mLUyH3GU4J3Vzew5vRACVjlPXerRlEtp50c9ztcq0gDCneqoowfXhEsaIjgotBJC0lAKG9U
fzCPsFXkD/ErFtZHNg+PjA8RMLdep2LnpgKEBErRIrikcvRO5qeKV5NQXBDBR5qdOq5IAjlHHylk
AUKVehybSl8hVj7Ehv1//bVyY0+bW5xBLgDamCxLdYalVUPkZ02734mqnLwkOnCzO/Fo0CWri1AM
tpJLf0XzIbHMfRigp/uD3N1co37o9zr3W32+RUJEwrruzzvOc9g8jz/7X49fpxOUX33vnM1KfERa
7tq0GWYoTANEEoEu0xNaPC4A5Icdg3Nr60oz6lF55t6OhuEh/R0T974Jo/ayHDlfmcZgjaFr8NVV
hmh1gJQ4TfiAd4FyxqZDnpT70Vd5XLgZ/IDocCFfrHoBMu7QzFo6CYGSud/ORYT8F2MlSVdjQAjs
M9sa/8EvvhkAJQmd3kTrOfTE98izydgthGP/iDd77PzaPmnCKk1d6vb2vlupAP9Xx38KJcqJZz6v
4vf1UW/lNrtiTjEKnPBSW91I/ulLJj5yDjH7Uw3abPDg1q+Wt4aJq56PGtbWZsGiZYbTeyI2toNe
vMF8bCl4rsp7NX7fXkPWZfVjkSKQcApCCUTuWzQf9CX9M1m7yqjRqe0bvJv7kO/MZHGhiunlJ+5P
lszg9PboeaTetVpOovGGyKtW7rUmaQBKiYkxnf1Kt2SFKaH6ZYxFwtGGH8xxpLGqx8ZESnvlXEwN
x4MsnjSElC/xYw+0A0bJydll2J62s9NlfW5osrqe75qii8Fhzp8T7Zk8i6Byda0J3e5BB0ab7rrQ
2ajNEGUjs+weopRuEEWhjqT106/zql8m8miXnr9D4uvEnUXrtDQwPsWCNWI5OHI2kC/IvMxgTKoF
H6uvq4k+0q0tctWJVe8NOSTFQRsBHa4t0q0MCOdhBn2xBk49dbXIXj1GPuQvZuwtU8g1hsOEYgKH
6oYUWekj32qZGUyRp64fQTbLKNCE9HuWi1m1maNoHoqSHXV93TKllRYccsgCtoNnw5azhVl9lHgT
Z8mpPASLmDCizUj3h4W18PCVajZTOGjwUuboHpdUAeAspbsLWit8DPGHC3IvA/8FJ6R0oAUd+q6G
c7OU7qPqXg2Hj2DUO50pCU6YO3VcQ7WDpzvkaOJuf+4LpP3hWtuMtwGBOinsibVRTXbiuzfOhqOX
rXWyah3aOrFbbOb1IZcahWqIEI1roUZZe0FylE1MCu2feyZCnAN/7GHt2jAit79avXYM+nj7sHjL
fy7s8TOGmn2mcV40KzwNWt9QF2Sql/IOBT6eTD58qHVi50JK26rZGz4Pc+ianmbjDkZWrlKeBzGN
vx/ctIC8clhZSScA19L9oPr2zz9TehFf8Z1VX8jHSUOITEPQ6BF+V5wdMbNPOw4g6ntVBOLnnV3Z
ZQTFhAtho9NIzMZKw3xLvHOiT0oEP2x2Prcn0dstHdp3Pu4K/GfUGOnSxemT3+8Tv+HAxjfoIz/7
zp01fmjE8FVqisQDnnRH5J9KZYW3lXSNv5K6QMFbNr16BLbrCtTLi/rswtKFLOnT9PUN+B1LeyyL
RrZZ9K3dXVji2SWs5TXlom0/uyzJGpmX9zm/ga70fYisDxwrfNdpeZvpNb/svcBKLEs4QyxlJ48S
eQ/ZZDs/pSYdmj0UcftXPutZw1Vu/813FJyEZum3bzXienlQh+JByj8cojpnaLCAbgyb7iIqZ/JX
UMa5lLKss0VJ/dZhIhWwwwsJQ6nZxxRtkOoMadGlmbzZ+upZP7ulCc/u0onqk7d61IkghCCdglF2
miKFfww4tPdqeYTiilamIivkUVo5L7u5Tc6pHpahOPwvcC4Czj22LP7Ql7FHd6QDmpet3Rm0d3HE
nhjkNqpB0qLqVjTZSGyLuDgAnZIPlEauixzxbvDiXPtX3nXgnYlLbVXqzaFJBcLai7bmcnSY5G6m
0Qw+gJGejilZB+8Io7eLmsMBmTB/bDyOKjb4daGZvLmibbomZvI3MOIjrGEGH/PqciUWPeYI/7KW
IuVf0+/JIRte7bDUpZGmN2PGhTtKSqWDeeL9+Hc8BSUsY0C9KqcfF7VePpwCL/TS0FVBB42QtP/3
o/lovh8Ub64xKiYYit6u9WtDKY4C6YEStxsJ0Uueaj9SPsfgdfRJ03D6TlJJibTwqlJ/7Kt+U1hC
BgvI8cL6xknF/g69cBVObBg2WrPtT0neN2pZeW0R/K/v47XCraV2FRkT1MgpQPriRAfUNyw/bB3L
bHhrd0mLA9OkWlYcp2Rng73HB+ZlwtsQ2ifwFRz70i5ozVyHxfVrFNUS5iccVaumfaYOOwTFlBjq
dplJve7GvoNmeRmeaA6XaoXjQRcPPwQHpcH52PDNOFkEzUtqLqbE4oIt6VHikY2YvwuxKaXTlnrj
I9N1r2rBkn2Pe1Mqf6KySMazi8xIxTRiQ6EY3LHAPikbiCTXzDPZdEXdjlJKlzxFn9ZHqaBrPC0l
ej6MKDKjKmCj5LEJZMsgVTeh7UgGZUBzRClEdxGBo4teq+j7VJK3Xfm334WHcKHfT2qlLgqZMAWf
ewfXmDnmVEHpv1HUqmHwU6Ai4TGLnzSkpC0Eyuc8YpluBAhgwiXpcRDQ8aZYalTUCf9fsYzO9Bz8
4KQ0Eb8uJ1SCLectW1DcPHpFwBs0GMTfWtYer2jpr7VBiv7pmJ5rDGcE05ywOtAEZp/uL37GrD6X
fBkLkBqCXBoTJ5/FN9FmotMKNAvhaBnWb7GFN7ZdZoc5sDXTdVKS2BGb9cGuV0lLh5Gc3Q1cLFvd
w1wy8SmWKDeAP3LTkh4B0UD1VW3uatB2Y+yh9/9N6lC7rA1AFxocvC6EZAmHP5zSTf6hxVLjzigZ
ylX5CQ1S1e+z/c5cK5fXFqtlNSH6f7o2Ztw8KPylqpjyLQozxetUF0XtOLkCiSvFRR9uYldQk7Tg
gxondHbTwhqtU2sGY2ejCIzD/zG8wVxOZ8zwP6RpIHxehPGC0TEjaXr3rTO9zRk4V6IH9qtHoE/p
XOaOAJN4nRLxwQaE9xro2E54carMmE8UuxmpDONUne39AXhBNZ8WHC9Ps4ONWggE3HwARaqI884M
/Gm/NsO+Lv94k3kPEIGJ/ddFmZOEzDlqWxgOStP8rTw+I4M8ZGTX5NQwIux9Lz2LQcoTTQyMpv1D
gSHHgEOfrYzA0RQ/N1RjUmhfW8ySV1RonNcU6ax2O4lA1HugIaHqGe8T0lHtYTRoHgSewWuCTOrW
kL9S6qAWHDdVYv4j1+gxNKrbArPuJvARo7vhCzANHeP+6BIAFf4bIUmVg96XOYzw9JZXn01/YKmZ
YiRVgY5hK7Eq/zWABI1XT4ev5aZPIZwAYonyp+tYPqVT88iaMeVdve2Ja4gNRGyGkujjzNWSD5jA
5OPKS+C/jHe+YHlVZvKCjWeBdFu7lzVxZ2/5OdE1S9aA3bFlK4gNS8jno4YNF6wWnFH+UPVRBFWw
BH8R+jkOhpqw0Lk5JT8A8Z5TLOluqkqrfpB6G2syZI7NFGB7HVmDbkTRgfWcQoxaDdwDv1jwjJUZ
RTXnXkNEQRIT92FfbKcTWA7J8HMcKOIlnY+j6ibZmmpA2Gai7eqq7FrghUNjsQYnr6AhAGowCy/2
9FQzgK/uqaGORWrPJtx8TN6OcM6vkAsCWNsqG83ZnGtTkbDF1j3c541gLXb6NW45GyQ+2ryEejfa
LMq8DKO5Xjd+1YJ2R6zZdMb9kTc2m+5IVx1fzJOBUdX0MyWhDzxWveV4kEVr12cNg9asQoMjXy38
CfvSVfKLCtdSvR0Ik+piEXSV32JWiTEX0VTPXelqU3nU+RO6WvpQz+dmqxIm5+h9RoPO8ckBONG5
wcssBpg8kV3MGzUuVe2m2tweDhc7pVoX2F7VHRMBBaa7WkQIDp7RW/0rnbHAM0E9Wxnp4dVFvLyz
cd/P4BweXouXb+gjLGHQkcLmQze1wETkJYThCKIVfnUflTCF5th3IaCVtNdaiumNlKaemmgo7cRI
dFL7eSGFFSm2tr0pWyjG8la247WY2SxBSVnhLYFpBDi3+bUznwDNTrY8tIvb8Mst38gWo6uGpLmI
F0Z5DO6LQMbVPwbY0eP/1/kSYAwxKBIP2dHd/AHU4u+duZPoBGGQySrcWHw3kPkU/I5iv6DRP09t
QHUUhkgX9PPYzzLqOUV0CT3MWYdfF/KcEkM53RE5diWy+Dl9oY/W9MHt1/jmpg3DnTtjVVfnYpmV
xF2bjO0MR23m17DeYhvC3tw0t0R5Ohm32aMOQ17PyB2r4wA+HKqDLjxaAhO7bS/Qs/nNCox5AQoI
MIr2rno64al6l+WD+RdYG74YfxAbWhNCahoaBmR1c9xylPnjToNNAieAf1ylt6EJm7f8KRlYNhni
3S2ufYK1U5BUYmmcogML0kMKrF/Dk+qjP5QLx93P/GTcDLkJbdPJO6OviIiRTQ0i7O9tqLKI82HP
64+n/v5zU2VoE8ow19Q+fyEunjuXNzC1MKIjh2fUFtJIYqedR/i8RWYdUR+wwG/VKt+um3nPZeZA
hLjZwQSdtdb+CaD/SoybbNiG3aHzp0Nfko5eOaMSn0WokCK+Bay9rtVE2BMDmIR2lD7+tnenoWEs
QhRnWUUztfjjVGmkB8mCfopZs7Fr5Y+UUGemiCB7yvWHcO2QIUX2PQ1ehx4IU1/1CFkVscRkFJFs
E/0pG14nuZakB3LO3ubMPc5PtlqB9ps7yfDMi0oRWFk51qinK8MgauygS7BHZWStRR/G8eRcb9TS
oB4nYVs2KBIOZ3IMT3433aGkMwQFA28vj+PXUkPLp5pvWkT+YVt15VVxN9g6VorBYS5Np4MWm0Y8
V/oe7yoTDDYxQMq7cxmF+B7u6oGiQxk7SWkes2ybecyqUyvZZLyy7GTvPkN+lKMmNVJcU4mvIwL5
WXvWPnbASZr8Mxd429mh8edjKmk/UkTIbVT0gfVneBFUAN7RdKDXnUPrUQmDSl6LPevf5/1KNMpY
OkU5wZGjgZoqPfchgKcth4/Kr5TgKIDjrTv4cd8WdBoreaPbbnDltx7WeaPEAhQsUTeWQHeo4Y2b
T9ofiAc+PRuIcZWrG0X6QBeg5oDZbMPKawWsq9+chanbj1Iz89gSoSLosBYuTzh7hziQMSz/OcE4
POrBqKI9w6bujB65zszfGuYNLkASHLbZ9Lh2bft3PoCOIudtGchx/e47btpG/mDocSeUsWejmAtY
TtePv1stRnZL73w8GjWQ9LLwTxMv1uNbvBXVmThUC66kuoSoH6xi7NmB3HDPVTrYAtxDQmRa2ZfA
h4NA0eCDVSJoD69kuPjo/n4VTRZucc4dX+SoVbEn/H2C0V6ZH27z0ccNyNvhR+n5tlWg2XfoSpGj
BpFwflh5d/+VvSUyOY6jKpZo6LDsbMIGtjMYdz7b88dp098aixZkpDWqgZJ9NWu69h1vnwsqjJv2
dR3jnO2Sb6CbVA0FTASxfssL+KGicHhfBKNAqqQ82tC3idrjHSVZkFI80BbW8J3LfWXaCbUBnWUe
ZT5sKqIeavS1UerdL2JrodWzjzKh6SWf6UqqCpROs87O/Ealu8YllDtgTgThTdsVezLGbhq0ZujF
CKUjftnsucjXTd+IQu1nHp6J9UQT3lril3adM/ix89r5No6CFdNHb0Lvivuz9hV5Nr6NAI5vIF62
10gKuQlZJljjRhnewNqMmvblAm5CWZtoMH3KqijWJ15GlA26CnVnXoH3Enf7ZtER99e9yz25oJJ+
QRInmZBUzE8BKIDGF78/IYzc1wXqL4FZb42G7qecnmbJrFjN77SJNTE5ey1qGVu8IQZWnCjNYvE7
FMbVNG91kwJ9+vXZT3ll4pwK2kB2785JuTHH36bOCkiAg496J2ZVuEoOVhZCB26alGc4d8kz016V
38rBAuJD/MuHAd3s4rxO5aKG6t+0Do/9C0zhKzCSH3oQo+g2mQM7e44e2+whLK8YwlehtMrKNz0J
z9AJRqm3k/RVgLegurVvxl0JUWGsHjAlnmgtSDQt+b9bt9VuvOOX8PYETeh1w/eWjj4v3jV/qsQA
BrbHhWFPr/udZgmU9gEnWiG/mL/gwodO+SiUoXGzT7jCSoabRAFj84/R82kry8FnDgICTrYHWEpM
6OJZKN1UWR0Yxdol/OaH0BT/FG8EbxDpNdbtBhRWNzcCBqOwWVqlN7QLIIQwR9KGVlYJXyxZ6371
JsXOCf/o7DkBXa2VLeHn2mcf/i+Iu8TOuHE92oGNPlGugiUD6/hkBH0+X0XAXAV1+PE63JrRVeBD
EmlLb1zdcAZesGdKpROfO5liSCZOcfG7FMVNBVckqk9WK8Ub3+TJ1RgiDujrHFIQ/qc4bSf0hL59
sP+nrcgD9XmEUA2oCHZdIa9V0iDKGUVyrZSJqESk7kjjhJsEvL1WzBS8McB8a9HXxdpY5ezO8cX+
AoxJQ+D32BqpxXeYlJvK3P0Mda3FByQEhMXJwpv4KhDEKxb4prev4k7w6t7+xjt5ONBCsSBuie9p
VTE8P6Eg24zakVDzQS7k6q0A0mfdDaEB1y9H7TvkOridfultuK3bh6LOlKqjjkeKc9hH2mGTjJ5l
0Dy/xgisczfhn/36zj4/eGfKr9cf7Ow6WDoPo03urxQre8fAFYqnVH4I4kh2+7MQ/QsBoxaiiC1X
eNTXjrteirH6oac75cuCOQE4Xz8rl/zNIU0xv3PXhNA2BGAMZHf+NfcHmoMr6ybD13QEiKYcRvhg
76DvQVPHTQ7rMXjCRM3Mta1Q2T8+sncRofZJyDXq0rdTqNYmdhkNUpp9UY0c1kjcXkyrs20PZTma
wsMAo9+Cr88hSKd3mxBIVPlnuZ9rTuv/t0x+tDedpzxW6YpneuM5NfzvW0e0S6LK7cy7fW5U7cOb
uNP2pTlRvmavG+5D4GSEBSGdLSertjObkOKEOW6kS41i5a0upSKr3IGeSmo4OjzRV186NxSJccXQ
rgE7uLurw2+XTqTlWFM4WP/lb5mHvkNzO/1HHlDMliubYGdAzo0I134J+Hlx9FLb5txO1/NOM2iE
0wmpw3Bl+XgO3FvviGPrNLYvCWTfZlhJZ0Tu1kGeFS9vcdkWvASuFjBMAYxl6aunn+Ru6WPBdbpk
D2F6VVKdSpmlQSiqx0uxoiaga8ldf9iGkSUIyZ0lky/bkcP3UnCQnVWT6FSuoGdUTyQPidlmPzHB
LzMdk8Y+Qk+2HbSzyFb3ioWKxgswbDYNl95BKVbCRj0SW4Uh+mTuRR5a9wgZvsqy4REBq+sdvgGf
v5+ehjxM7uDnvtjIJxHhZbuka9YTUwbA4812RpUiglbHBERiQWNB8INwhtebLWKsx7pP/SG1xz3d
ySuzD7x5Pt/IZrP3JP+4GuJ2fVN9c8QgLDWaQDfC/R6KetYjW9LmoccOYbyEEAJwH3rsXDQODlWO
f7JvxrUFIggWnaW3eeQTjfpE438UNsNqkmIaocjEXcgR08eoq8nRfbgBRm+NeDBr+lG0Qzac02Iv
+NmqTCpeXsf6G0mknHJUGltXSetueDcqGv8ZxdTXzWZc9USJTWJ10R6jhBWu1+EAKYWBDFCppPzo
whulSSg0OSxzzhUnSKtGxYzSOFbljFDz+KHwYOjtlXsIOurZ28rfibCw/L/QoSKekpH7NejruNAT
lKuKEPCjT9PwdGmEWlfatGWI8H8DyogM73P/o+AEY4X/0DjjX4d4yaWzhognAR2S6UQJ3fdTf2zv
KXeXKW4a6ibk/CRk4UXvyK/UwVbqMBgrqekesFGkusWrXsjrkLBLyrvOzPHZm/cFI9YFiHTc0TGM
qxwCAOOoTtXuuDPS4onJ69oyG75FrS++6dACl9C2QcALDXO2j/yOjG4xu9/wWNi8oCniuL50iHHm
vyEZthsr/f+K7dkMsFMX5x6zAQzNaOEkXppKwEqClvR8jptS7wvQrbvPaRSDKFGf75fAvsjwfLIB
cA55qL2oLKEn9oU+PIPqrUHqyW7l7M0m3veuHn5gBAJLQMd5uti0OwUCzHgAnMUydKXaoaBkyqdk
4o+y04lATqvcSPd+ROrz+xwnXN2ibLhbqcUrH7u0fMbk1gtCP9nSHNGvj7T6ULHb0REAVfj5LJyh
cBOqjE9U1QBGv0nuRm+tnH8AfFCbKOxcEukzrDvuU1Ww8xQzZ5vh7CQC5CW2GeTyeimoNKKPPGJj
QXEcH3kOzOtd1xDK0veYUyyqqOCFoYItz/IZXr3DA5uGREKq9FS8YQsxNoG8zqaqVCLoO+6sb9fP
kWPR8143bgf9eXfDaUtsiRJo6VmjvbCENCDtuckOChSJoSU/d4SbAJwLxSeWEa5oaXmMeQREG0BB
AZnnUY6fREOMKx2Jfu3mNheH4WjPkZzOWHadfL8tTzP6XVaOrpheHvvkXAMBOLNn9MHGqOFdEvir
hDuVVVg0elYO4B+6E/+fQIp/Jxx0t3mlRCTv1WYymsmNkCq8Ij/uP5S4hxmc3t+NThSvvCTEcQdg
iJ2FtFdwFYR8msLJJSLlEDn6Y3PxQhz9uUNQUhEnB4cWf/J5VCBBCd47Wl7vbwehvmBcn6uM4WqO
dZOhBPjautMDo8ZDB7GJkmNTCl0W+vF92D/h2Q+TFNSEVqlcw9t7uRum+9MGkGW38JCIc+4KLIT0
tmPzlQy9AfqyS4PlXc0GYioc1QMs0NWD1IrJuvhHIrbUDaLmqqyZH/uYBsmBm5o6lovE8DF0pBpR
vcSu9xqa8eiQtNJZiSW+814RYDGJmXhCLSIDgtrSHAgJ7trzxDiTfDcwNKGlH8dRKhri9bVleupx
2SjzIi3n7PU7+MfuZqENhLDO+TcPWOoLDkDHSZ+l5uBt6gZR1f0uRRXa6ERqUKKrFWMpyhJAR56T
LsRC1bIZemu6kc1Kv7QHRXZbcS92H79yriJFDpylhOgwV0uC8gcnTsKfzkcuvGZrAv3fXr0FcDkx
Vy4Y2DnpnmUkqB79SvWf7/mUZLSBjp1FylHLi3O2/O4qoH1vxTZqV11Kno9ZBGoBEpsPdl8BRCK/
ZPVjMnFLzfF3yIDoGFUeqZcybqeRQRFx/7ffnDTXZtnUihpffnG5gojlI7Sd+iJnAjCeFxmpaThY
vB7UzZVWAc9uBYd5h8V0E1Hu1K4JjuEzaaYnw/S7+CSDL2SZlE5zT9xhwqZi/rWE3i7LevoKWm7x
dDXjib7/t+w0UMommRs59CuXSTT2iaMMFbUiZFVTxcfip4lXgC7266fbNq+pmsT9xNZvi9d1q+Pp
OB21dl2+Bw+WL95PNfne0iC/xkgvPhtMfKcHa7g4uOYajPQerdKoH0QJcdvy6iBZEt419dyqVJG9
HmU8uuKeCKla3jwK66OHREtdRB5XO21/ZiMF1uuZ70n8kyzD/UG5xYXhR2OGYaduFdhiBWMm6MFv
hftoUONF0+Bz9dl4Bc3Mytw5UbYuD6dsT7GFfLCniLMYCjEZEs/eqtYT2RNKEakq0+HP1QZvTKL6
chRxgmJwxAqH2OcC7h78eyjGx+27u0fbhFGo1TSIcoTzu1N6zTlQ1P1Qt70UBI9ZA0AYbCROgyA2
tELI1sdOoM4Qo9vRxwRduwGRbYysMdvGB6Sdw8mlMd4DwUXxxsBM+XtC47clzgRX9pZqNBqh9E1C
AfGDExtExw/VZvklVesecx9bX0VeT62J3pSoCJKaSeYYQD4PCjLaoF69U6H0k5tuN5XpqKVZgJk1
Mlvh/iuAOZ2fHwS6FJie7vbSb9r/aJaBes38ar91WyNSK0ZySQSN0Cym4l7UBvCnn/V7ELddZCHm
hEaiVU5zUMqpBXHiNVaWWUmNIRCC8wbN8z9x2JerSe7lOyVRVal2v8CxK5WZoDOnzo2k5ItF83Xf
t4bnlAsD5lTRP16u0Hzq3kB0F7s0tGaQHIf+VRWW1suQ5mQpAiEcSoh+z+Xh8jyxUCiwz+qJ4l2H
OuTTSRoEFE9blx87heQki9Afi9aiCALwHn7voa4kydW0pnq122VfCwhcAPDpWpCZ3FEMSDTHjDXD
MK6SexmyaVpQDUI1wjqyt6NCC0D78Pp7Kv//R2iy+pmjcrXYDN1MFuxLNgYrCOhQ7kjhd94Fsh3m
KpqSKU1LxSqqr2HtaSXeL2hQpGGTGDoX3ShQ04hT/1qCSlKvgRgvvYypK78+ia8Us2MQQhGwL9XP
N7SrF7VriqWhNeR0LWBCR1dqBjsaKOVVlwu6w8W0rPOkgfKViKT5wudyz6qLWoeNI4aGmuWeNroH
4e82Jk1y/vk6ooOX9iDhz4otaZt5RZkxG23lH7nqgaNSrEES57kJhtO8Ge06f3S/zISSMFvUpbNE
t0kUtOhJUwQm747X3brU8dCeYzIPtxzF4/p8JPpnTp5vn3j32sU69atnfzdUYvn7nU9C1O4Co6Kn
9vmUPCEL953KlERXWeSrLV2sbzUM2h2FU9E2TneGtw9gV2+SwDmH6gXvRqiKXcXgczIU5YyCWhDQ
i7nf/UI3mladV7NKZ8xej5Eec7hl8Y+5BaimVaOBn49fhJUWx9TU0iGwrkj3aNIKtrQ2xFkXP3To
rdNzJy6jmbL0AGowvJm9fNt5+N7ujchSzNUemq6vVklkODEoMyKwta5kUsKZtptz2vA1WXIgyz1F
0Ri9b1S1UH2lFMdQmHD/4tC19ho+OFf03PK+T6UvWmc14Tu7jbZx6LOg2QhmCFGq8YHiQuMRiila
4xklprvnqXbQkWulMNJNEI5QCb/SaG90xRMbTx3uo64J/H1QNPxWKDDezZ41gUrQBa9n263SCCBJ
5FFhtD75MDOhZW1UzvSB8Bon8uhHZhZLMoogtokId10JpC5iBsvjzPoMC1e6EXJ4exLlukaFOqW/
NqfKNMflkJRX8svorBWeMCLEhaQfAFeAqIfG17b5TYKCmFxbPV7ldPawd0HRMvH8HF6Itrro86Cm
IIUL9Z8/Zrj5hjw1j3f/O5zILpo/AastnW9oq9SeWpvtqSsdO1Z6PdTAfPQnx1AB69VuAW5PgD4T
OtHT/vZ9uKFsBK0dW0MAOb/EUTn3Yo0X6fjVW8BDK8qBJqAt5MA2xPj+8pQIYEbTkvKrG78c+p/p
gLJQtDYpIJkxqSg/6rXFGl5Igp0GRfdm+39B6rkMS7ovEtHss7oxp4t4xR/p03Mnw6w3alDKE5Vc
KkecI5QxqeRFFzIod9gg+B1R4O1BOHxhthHvIkezcDdjR7fgPQSKizxjchOkxijV+Jf5Cd9c4yNm
iBjs63ULTPvyY9RrxuRZBRDRxj9aA8fh26WkaXksyHfZBOdBHtBGNH93xZNN5gRWanBZXZFX+ARP
ULDfqE7B/lodoBeeEUzIrk4O2J77+b0bUK+9nHJJXjiY5KYQrT+KeHbhs7cpIzzyafYmOAfhP/GS
92DrTlcZGojrm6xvq5cAyeQgpePA7liF+aITl2rsDIVkigbTqble0RrHSV6ccnyg2gMdXkk1nfrJ
Ws/fUMypp6M6b2z5fuUPiw7ld0Rf16SofLBMTs6t5CJwYcsCGpbOZknCTrYn3/49I37zZ4ru7eLy
6dus0VWuaQZmRxVA3OjCWiY6okTx7NBD+80j3BlH5eulH3e52Kc9A0RmO/78T+DE0aQyyBXUWgOW
SfJLZElJWlHyOxkz5b/Kov51dkpmPptNNMqSFUXDj1NyUYiD0zXHdYwz21RSsO+reeQpwbgI65Wg
22GVJDRcv2alPYjGy2c6QAQ3dBR8B2IP9oBcZH43x5qSH7446mRyJv2w86eh0ToUXfFCPLYpUiZd
D6FGsvpu0lTicyaQ3fdjRP/wbZoKxd3RjpVCIpS9wmZrCSIvK+QX3MDyG3fY4r4omEwWh4MVbehv
nDdS2KxwfB2dCg5Nt425wLmtIwS+r11NIwoRSHYQHrIdiXKPialZYtMnCT4Ii3CPzIvUbpgrL5UT
0Rc5llqXzLgOLZnSl1lCHpPzJFbpVDRpuvdyIeRf50596snsFVXEXA/5oC1loEAmKnvuZlELb2iO
HnZxBrVBPWABBU/hiUBmY68j2LqTCOPZUcsILfF+F53hBdJ8zgrHvyvb4jnakfbUoeqTNGUjM9hp
QVPxZ0jIQAu+KNLa1l/4SHl9sj7rkkTK/hzuVwhI3oS70s2XaxaZGf/Dh5AOZf4AXnu/eoOYMBR6
PYGxLGsjnP68ClRLzoGjcb4xchHj4Ca6mlj8w+J8xbU4fQ9b33qX09rtmXmYDsgrEv5m4jkkLJmC
RdIsA2lwsrjFX8NXWJweMvPff1NJNEpod8REL9Ta8MTOuYPANYmPaZz4MFDSLu81zBKP+HB1Ilrx
40hz1//w77KQtD7ynRkvs1Ja6+9x/G19B9Jxyu9XI++sEBkV4qXG+7YFnd2OL5/nHqEtbA2rWucX
bYh1caKW7EOP6baBwAw/2CHdzNEv0DU4Zu7Z6/+hNME/BAK7tFGPS5Jfv1SBlSE6nylZ8FTWaBlx
sYTUu4KcZkTygERIMhrb0pc+ejiqW17KnLhLh/qI6O1SbPOb0CUIRwhydHqN1E7eflKjEgWG+R+a
Hz7TEMeRlnwzp8CL9JTpK2qZZbOp/At9xZqOzz0/h8Xj7EWIa/kObqwjhIw6r+cs+X24xthg/1Ni
qgq/VncWzac0U25yQfDOpCY/dHC8JwvmZtblPJZI/Cn3tW1l5ZUA9W6y8EMq/GcX6VM1gyUn2iB3
/Npi22LHCfh9Bzaf+AwKeuyh9toycP9vaVXXizctafOCZ6UnyP4/scfcr+ZjR2MqFE1YQb7soFCP
FiYrrW9lmENpJZALTQOOSZCzjOS7TVxGKG0X2Qnl1XZQb+uIVCaDJafhwyHrJO5X97bEeBlpuShg
o03jO3DXEuzqxDN9jBipJd9Fij67VmDbYTUv7sPWf3Fr6J61vKCwYrClR1hjzGi8MPUXudxH6fEd
CDESVh5qEsYygW66vYUkxdImXFGThTiVTzSRZtOtecCnFHRbv+m1kbNaVnF8HPhnSBJCAwYVa03d
GqIgB7mNMin7DlEsAOv30GUKlbHT+0gxYI5fyj4gKY06+0GkhZZPFCZ7VSkx7Lnaam+I6ZXUC6TN
6HeHKTQT8fk+bdjDr3uJxyZYIhg8r1KVOTN3vRfFUtRAB8P6fg9MmarWzINbCheicz/8S91cptHx
DlAB+KCW6FA4BK1HODGaYNwPOKTrdufZMZsfCV315IIo0rAhUUZSIzF5FKfHI0t5b7a2bahODMmd
UqrbkuglqxsJD4IdjJ9/d/x4CZCstKjTq/P8YrwyXgvQOG6mF7VYfQiMTuHGS94o9SeaD6Oc/yaJ
ORuNvty87gsulITJl4GlNfHLCdzgQP154JzLaZ3udSBqBsFrBFiGJ5KDonA3tIGD8Ebdxw718xiu
NTX3o5oE2KCL3EcxhkMerckLq5ACJIWzf+ImGx53Pr6ZGrL7MGsGOebWCqAtpkNInxBysDQTKiKe
+kP83dKObpzI9kfh7x6EhFGrFEZ0w4FeO0BeEDz9s7SSenTcewNK9mBDE6L+d0SO4bah9ZvSxiun
ex+CaWbWaRFK0OD3pyUa6bvUJ1AYGzz6VAi9h601N8u4H++8KQzxwGnMVnm8BU4ONR/7qZe1ibSa
lpsAZoHNY2bNw01W5JrQ4kbRSnQs0Og/Mu2qXa5/BHF4XdBzZ7z10utTkTnfmyPc0Xi82jeTNa3n
jdNHL2Zkc1y1H99Q19Ws8QA8cXJbBu2nI7GJgTvCYE6FRVXRwgVu2DeivzLaY+WoonsXr20EW382
zFB+x80MVx98qc+AWjLffbmC30gpp9uZyqu97tp/D6961QDRG87HzmgefNkSiXtSW8TXfc95hzke
UDVt+ftMVrCGqfTpQDb2UonxAVC3cnXUmUhZT+HVkIc3Mr8uyu9FRD7pqb2BTAaCRqBirzcwWk/b
rhqWp3fgPm6mQ02KGrWR4R8FYE3fcZ2AC6c5XD8WAJRk4NOuFYobUrxaCuvpHXCQO0v3jdi68Vvi
eXSMaBAyGTEK04Q3PMrJduZXZWNIHw0XSdne9RpXpK7/6Jq4kjYoBltU4UMM0LiFTlnMkYFuu95O
d7JskSq7R+jU5vig44VMP1ajgBpfdZ4fyKTIICneeEP5Qhryd3xWogCYaoXsa3iWd7RKfLAaKUqB
BsH+1RWBPIZgoNQMZJd+Kg8Q3fFchSeW5LNvu67ACIr1pJAsHgxgtIN1SONFm5VdS3ew07mvmhyI
lBZCkUUc3PB7hVof9npppBWzDi6+yt2RE/F2+CN33r3YV5eP/rwMBsAHxMvOznWHKuMJ/L5KEinZ
O3Xdickrhp2vN5BwFw+QmK+0nVcl1qlvyCb0LgYKy8B8IYffG/K55z6favMgPDRKSa+owkRVwz+8
XR/13Dm/kwXnAByW5EYheA6AuyKg2561hbxH2VHOKE1RlFe1P/7Gw0r+Eefm8D60mmqL2kTaQ9rg
1TiELJiNLT+aHTUCAN5cxoFTKRitzKvJ9ZYfYr8WVGTuJFsIsY7i+BsuqyZJWO2wbDSHkzADR0SF
61j9EdCBzjXLGcgCgrJ/ojX+0P6pyQJ/1tfV/kjMs2ITsA7q8PvErytTP065PVDRjaJkPbxw557L
3iRBJcjeS+/r6X8Cka37rGQRYX8V5aLQiD9CjC7yjJml1sWyRncUAM+u273YbusIbnfE0O29ccRF
S3L43ZyD4cFsOY6SBbADX/b8gpSBDmYUCRFmreOF29sOfIOnMz82l3V1c76M1C3WnLJnmUg4fnU5
CTssYLRSnDIyL96GJI26s24GpcOHCwglylp1wBl+Z47e98i2vhAgsTK1tWmjPEhJUiHYC/gqxok9
PuvtHZzi5RShlDysUj3/HZbrtFCxlRpVnIE8Ebvg/99QTUfdKEzgp+STSQFA6Sods+q8N8LwEEfk
sw5z41TPDsP3eWHAZbphU+WOw2GtMn2Y7cZvp4E5kPf96R73fpYTrOS0gxuNEBBEg1R/MbZvkETS
mXCipGjNQsCqIGsS0TFIqhr4tRtQWayvEZ9tPgrcGQ5hs212QuAIYPZMduDIH21FGeWXA+ySE339
Q7B0BWeyxLeAeabDgmQQIDYCDJ39lUxkxe34jap6u/+NDnSILaHn7Yi/OmGR/GA2Y9UWhfcQgvUt
9F33volwId04SXL/7fYW5FKuns/dUUFYDGRMfUHJGFRy1XJ6woOnPcSW+xwBCU20J3mBWBQjpE7y
A7L0/TY/+wlDTfXEjZZC3MbmakhCXC4hA5vSgg0FJLwuHa5XJCBWHfsHiyqcNU3a49925BsYNa8y
NRbcuYib8pbURA9oTF5kIXXQNeTcyxaHbW3up3JUy+OnbcDBKqKzjPJNzKrEtwwqaxvExkXFjPmw
jko4+Q1nsrNrhFUfvPif/FLukjknRK1AdACVx4wp2kf+QhUFMvk5ifFExLQ4SVa8gSpNeqWrR1Ye
ty30GyeT8fxmpVDiQ5mrg6OmObwV9lNhCw2G9mreorUooYaVvkrFYwogAmz4NTLiRC/pDPT14dui
uysKjapE9NhZ9HUTGz7uKFlnEAZCL+Gwvy/5c1uYDurxa2vY/yJl756MbDbPDDSWid5vWpht+9Y+
Y+GLi85FtASQ6g7pk37zzxKDendtKgHU5Z1hpOmtTRHcDGxkaG1SeBbDVbuXbr1flOfFmlEPKw9B
kotgViZ34QJJkPIYJ8TxfTY1xo9Sox5kvDDLwqp1Rn3G0Qo41LYkfTXagaanA+zrVSrM/O2EJ9Hs
UKAQYpLnbVHEDoVfiYRckaXykXSTx4Ju2O+RQwEZ8oc6P7GpiVu2U9oomCU/w+zhN1gw356gpVZm
ApZIDvRKupTY37wsOvrOklEq18NDzzweI1kzSz2al3/Ulh/Bwc7FszVAQDVthyNFf2HTcSJUlej1
SECPmPl1X/X2SLh8cEqOmZHX9UDYtLAWyIzuH1UL5DiIhqXMtv4j4RbYRIL6u8I6kla+ESOv1c9Q
Gx4htmyLUUSlkykpuH+tNTN6M7Q+1+J1RFLWLwcqIiPpwH7eq7AMAODVD+00uBwIQkQHWaOmw3V7
PCg9fYrtYFtd0l8iLKpn1Fn5FaNfC016pIZaOWBmde8c0o1ZNLq7n1bCggyLqFNIp5wujerA+JB4
ApxKcZSvhfatDp8KIAZHB2qEkiuP4raVg8Vb/FVBQnPzVa7X51DeJGSbFqhEtSUDQ+p470MTXfZN
GGE6FEdSOLAyX9wPa173Hleoo7iluxbC4AvJHu7ozfAfs4tiRS/hr+CQGzv7QIH96bHSx8ZDOiAL
MXy7NlXGMHCfISYGonZW+N0qp0TnSZBt32juSVyY0MHuWRTngL/r1d5cKkm8ZAJUGWF4fOcvpWFY
cDARK9EivYKQgjLRn/0cBy1ZVcXfa8TLRf8+gPZa5KyRps2DFZWbnj/kF8U58bwlQIgzB0oKtSNt
CSJiIEzcQsM9B4JyN0i49UohVE0ZL+QL0YRVYBtRyhZ/DLdzu8IpXfaEpwdxZnBu3yDllXZtkojr
yK0xswDcg/m+PrH/75eYBWR0+ihl1DPz5MEBhAQcHuItGCtpId8cnQMvkImdR2KNP30hB5ojcxEo
2UCEQGVlvLTstM8fJ9Y1plbsv1FXTj2g3iNTqQ8g1lWKtWUWhqQboGYOE/9yKrCJ+MxCoxp6fRET
AjMI4FRzepVnOp4lUTioWF2aNjVgVfZY3MxszTbXdeS3FklzD+88fgKzgTqOGP1TqQR6JHW0k4l4
1IMSZ0PTuXl67zcRTAZ6A1zWdwCHLrLElBfj/AiuaqZf6HBb9j6gHdYYd4iOUp9SBhmT9gI+gY4j
ZhodWYGB2aonhAE7OBsiIJlpw/xPGTvm+n9AtDcX6DiH6z2zktC8Ip0yduveNoaSo4O5QpysUsYr
S6kepp+qen+vv281/rq3XsRgc+SpjylWGM6iSd7ObksYXDkmCpFVVamzZ1XvxPxrclVoKPtW3D8u
EVGaL+BwzfKcawr9wniykj10yVIySrqCqqxi0wm5ySZHjrNGzDMQcEsj0XDXk7P7Qtr8m0IA0/fj
cVFLlvN0jd8iwEa5QLdplpv/p6CYwec2FjWTzfhBljke9c389YFUFkRYjvM0PzjDN3dCkec9JRcG
sX0AvEOLkq/IVnMEnXo3YEMSDw4riFXSvo5VN1EZZZea/2hLFPTdjSNVR7BpwWV3ozqsetbU0bNA
e8pEXX9FM+EgiAO/3syhcv/u7E0nAPwpu0X/pnfoobQ7mWv67AcIHh8lxf9i+bgnGXnJksUWBy2z
AAE61IAiXcg653FIaKYF6pW+7gCgH3E+4VNFIDgLpKVai0gRasfqSSdr+o7g+64qlPDN+EpOcLWh
/95bfOarAnLaxhF923ciKU2GMlJ7OaIPIUjVUMOWQsMmRO4xkcbkQv+EkJOpR4lqmZMwFmC2UOz2
PsqnrTJsqjM4t/dGg6kw6jjhr3nimOnF+8UhmCUvCYMZw8bBu1Rkh2SiGk4veZVrwgTfwQA9A5Fl
DesxK1MBVYrDF/JzLgY2Vvb2LI3/oBnpmxzo2FzGE3u5/+YZHfXSHc+dyfwUcSHuGFSN0ZfRA/lL
DGWh7xqd7RT16m+tC2bj22mPCAjNQ3zb187gZYwi7+UsgLkSWHqz902YXrmaDi6svdp2y/g3J0HF
EDtkLIfcXilpbc8w7OmKQ4K/oSN8+Wbifl7KAzDtq7kSkuEj1NmzJR+MpArFHxYVr5WjhDSUogD+
rTUfG+7IPQp1NhnITpc3wm46rel72UN2kLNgDMIW6qZtwYxl1ePPSP5pZtuwFrWqFAomOxlngvHn
wtMHlWhGaEmrqWetF05zUGbQxa+4V/6djORQKgtqSK0yk/2zoAtQybAgKfTpsUrM543MY8u7PzNj
Cvz/brvQ+3K1p+bv+dxEb6+2sr8zUl1NEUUKf1QfA3+eyLYU2DoFYfCds23pDKm71TCEGhTjOxOK
Ka0e+5tbMYs6vg4zWwK29fUaTozHrhmIv5hUeOUt96MkatTVe+qJJSoez50kE83mLj5FSOhxdISY
qR0gQVYQ4Aidi9Cvo/xH2aryoLCKppjfk5DVq8hCxyF6HDAEq678g4iILcMeX3rttXQflruGUWQT
wpKUEZgzTqYMAb+I369dubDKQKgIr+97YDxoAiIokp130gfKZsYbd2i+8AdwTKxpXNm0Ez57s3n3
8o519sZIXHm6aqBn2HILtXp8eODCQLaaEeSjdwlXPt4Z1BqywBgwJqgVzYF6lRToRgzGe6e1xVhf
9m1JdVgxOf2c7sKuMBft41Dw9pCfJ5a1sRUZc6uaIqrkAOJ7kyiCs0H2ImCbBNOif7OHZLdD6Fz8
uU5GHhKGJdF7t6qpT+GZUelTrAfXp1HPj7gzQR6vJi2I5PhtyMIAMKC4Th42kopy4SVXH5f9wich
jJQdC98NNs3hKFsAo2OFX0f0Z6cyvYT3WMwgsd+01TQYAZ0R5jy3N0AxG2ybjvTsyz3DwFtCoD4y
l2etNYqXnFZ0nTdOHt9od+ldToCjTBarlFO8V322J/xQIJVO4kgeqxTKXLMam3PUPgT11cvS9w9X
G/ULAv+bNd0SkF4OPGS8hMOgIvjXPxCcSTDezRJ5Wy7LIbm8mGs0Wzr8XpmriMyxYEDh/Ijoer9N
xjzBoo9QkAYx4GmfUaKiiSMqV85CoJHkPIEzEFcoB4BL1A41AbNEBEus/p01KmzaLp6ps54i6Iok
nraFtNFUvV8gPTweeSpWji+fj/MJpzJCbQCWoRBb1GkBsb2uK21JZKTCv06HMvK1SORrOCdgXPU+
fGQNv7qgWFZCOE0dX0IeUKS5/ctLJvP83Nv6GhUgW7SO3LF+h8zOXM8foVmyd0CcKHOdcQ/O7hfV
3MCnjIMXoFMYL8qSXYEGIqoRtbO9A0asagatV0U9nqM2aQZu1JGpmL9wWE1Y9WpLwZHIwPW7V6qE
/Qd3wAYubgWbGoBUn0uAgTRNHJQBUIxniqeZL6O1wUyy8OxYKZ8plFEn68ID6ZoXcfMNZxOjR6pF
JIc292IyAX7KyxuJ7AcJrhIDTswDIMw7GqZbefqnuLunW5ldsj5l9xfyzsGhnr8vkd6vUL3Xl2hE
GivfuSzk3vH/8QDs0y4zoplocTwlyrRrxr9j1D1Q2goRSxN7pypbiaA2ycmi/RLG1PiuArkDuS9L
otkmZi9BM7tJrinSLluE8q91SwWhpPL6JOnP0PxScDtyX4DRt5ZlYes+TaN38q0BhzEw4Vi1MBJr
qqL28PsUIWSM9tLlWjSWCw7cEDm/IzWfn/ehf31TNr0ZlBAX2OeA+2oVcIY79HEklkOuCkwUlZ2i
7Au5uohluqMhsG0Vpq6TZ3cYlxXLnUVpe6UCK2jizQ1MxtLwEFz4Bg2izuTf5npGGr4k9LdjHTBE
691wm1yP050uk9HJynKDvH0GY7pQd6E4OmPtjVdAHcNKF1h7s9awzFywWQ8wPPONlJ8VAX7+0dKN
Y67m8LvaAOSVxR/hh2ezLTtOXzkQ4wvdlbw7y7XDzW4gJQW2BTtaMurdjT1U6OzkKAk2fDNevZp8
QkRQCy90lNExWK1kCxpi0i6oQC/bD33y2qXG9bWNwcKwXltW0Twnj3O+o3XL7vRnVrFfjn0IjA45
m9r2zLRWCQoi9PAGiu82zLhctH56eUFF+Ok0TKBP9rU2Wg5HONSZkigxzo/uGH0JG0a4afhez723
YSBfljDDj512zPjcKBUrOCiog4j0WmEaWV54Tj3JSeaAV1FI2oxs5v9jc698cGRk26djx4PysEQR
7yzHUnmI7KMwIa++Y+4wxFilHLvnNKauEz7/Tug22jEmQqqF5ho7bN3QbBc0Wi5r9GJ2eIz4ogIv
7iN0u33hkS+2OrnCwDNQOJMyk6VzMmWu76rmWXtVX8Sz7KWVJ2SAQMW6lqUQuLpuuQ3UU+W2h4Kh
CddhHcTNlySFoRdkoayETbfsGglBp68CoTKbGHMayg21sWiJ6FebCZI29pyT3EQ9BqX5wRlDiuR8
xEpHR6mmemu6UJOC6mxxFzZXl4NgKTCTqzIEX7yUbaCoDjqszlVW4595fGfnjPhtUhoxPe2NU4+q
0CHRfv2hGLivlGtLd7o+KMIbULpl1yc43IAAOcqOazrWCM2rKmkvLT0pksWber/qhqdKGijEQlui
13uEE/Xo8dk8eAF7cKxNH+5d4mieK2G5kANK/eolVL7m6AUWhN1DfqQ69Oa28wuTR0pYos6wJg5p
qx/gQdkChNDOrDmveGfW1rUSJhzYHQtjchJuPcz+9tqrokmw5bjPOSJJVDy+opkWpZZh9mD4KA6D
ELQ0HkaWgNcK4IgB0Cbx1sfixOBBLlBsURQjf++N8qmyJ1YLcQq75DNFZoCXOkteHbHarj8/YgG3
pmzi4uufZEdMi4ZmHW+ITFWaMHM1t4s5pUKXIddd81jQTwuAUvVlalSPi6PJwiDEUcJ1ULxrASJg
0fKBOECpl0BU5A7cHgIroOu0z5eQ8+0/dIWfRtPMblwWVutA5byTf9nRgpOK7F1eVfVv65X71xvV
tdZ54Z4zPwplGCzbc6RFKae739k7/0m6YSz6W5FrXE1kdGDKzSs0i4NGKZ6xScs+iqB5479Pm3XA
uEaUgGNP+JVgKNdbYv0udnBVl8yhgXIC8Acb+OUyesaybg0SuG/+MrygZkfgzO8zoAxThrrE5y7g
gvsRiWUgc5l5PQuQFuFRkHSNSEPjOVWy4OPxjz5pouDmMmVKjOjXxKFi6bj1r8P+Qd6U+2jYS1Qu
s5LLV0hEIpTnnj11gC4iCp38d0vSeGpJ2emZsKGH6zalCrygNw0Ekqo/ArfH5lIBzl/MIdGjjX2s
0sEovK7SulGwJrWm8TqbL4nI4WPji4P+Q99dHoBRsWOVrbnet0st4dKbBLr07xJtJrRzyxN0faV1
i5atNr348NzWBas/aKo/pIRseW8vKuBtgZTU420gLBbv1XNuaXj/d059KALMl9uWsyqeMxWE8RXm
hdTGwrfBNXMHiwb+4iJIOJXIt/2p4e3t7OSfMOUIsWqSIfuliETgkW23nKo0+Bs8O7n9rpYhRTBP
ttmzujRr1/J8b/UFxRA3Y3+kawxqPjg2oROaG+M71boq9Qqsot+3LuzPw/WHyE08hitkD1YSx7nu
I0P8Wa5Q6hUSlZoFhU3YRel+0PgLFw+zRfaZi4M9J4Err6vgG/8c8ssjFAYmByQD3OfRJb5hBToA
FnqotMDoIFKEehzFPON30Nb4UNeDnuK+I7N3MVOhC/wlzLxsSg6vM6OsU9j6TjHxPNdDI2BvNIRU
tq2EKSE3kIAH14spY9aYe36NnkdNbOa3arNhl4kAIgTC34fpNGGFgMhl89ZoyIdiXS2g7bxnHCOz
gpbuEOkHmMXpoBaz5ic1QjgzWve7+CSxLJJ0JlzyyiiVRorY9sB/+agTDZSD5hJNeEDJc8tphvWo
b98O+1DM0ic63sfHF63KPsWrt5IX6trwMkpmiq+D5O3E2qzENnKauxoXmEo5lvjt2bnkepJMjV/a
Uv6NSy/LTdpRKwx0W2iEGS+Oay/8qwdrBhf8R1D/xNhH0JRs6jTvqzJb++OcJumhRcz8E9Wd5zW+
RBSpV+e7f5Gel8JHTamc5rHPj6siswOPO6htIHSG0PvefKxNBwChsLwR7tjkmRjk6YFJPhUpvaVF
j8AXDF2gTs43jx6gQq7q0n+Zkl8joLTSa6PHSYePrrQ61As7Q062zWVxdIo42B/+r0B9k9KKqYoD
zMel7/z1aGLu2M6RFrPLCN69lV523fNLWbfqj/lD5guVC85vgMDkcww4cN6Y1De+/avSvspSrnhc
k7zbSDe1+YDachmi3ITYmDwqzJTg18XKAdDv46ZxxOaCTHoZ87qK7AyGZg3tAqCrVL+wV80oOI49
ztOSvmb3oo1dsr9TS9Lhi4pzGr6RwRRN/PwHbFoJc0sNfdRYLo2xa4aKwEi4AM2NEHMjeBZ3p6J+
zHZXJc1pr/MelS5gywBfUPx/y1Ij1KorHSireSDjCprZFHp5vBQb4DO/ZAN0z1uUTr90xRzhWiPx
Jb5oHR3Px44/j3i86ulWSKIKTtgqgU1ujL2qQUPOcptg2rVUUXq33ARjAwPpG4eQR4WGjur4WiET
3p0cTqK1fmAfTdQDAU97McLGyICnvR9nWA+tweutu+orr+sKmyveONwiZ4ONCJSCpCC3OCXWT8R6
auKSddsSQRbQ850JtE+ky0GOmsc2UjsMY8s1nd0ROKp3BM5VEH895P6nLq+62CD/uR9GDcN7+xpB
wqcLWkZO8xrg5Vmp6HqlbEY2zSQzUYvXgDUk3MauV4BjhRqdtp990sE79r0DL1V35o0XIULR6Ppk
aMFVyXUF9DRW2T7KYB688aKtXqIB6fAUGhA3+Cs3PCo5Y0Fxo9cimt7/l4qf87jfvPuk6cU5g7Vg
3/BSHXA+Ae2hDtVug9LMaBln03yYbe+XBXylD1E61pk8HhByFlRhxLPkBfUCdgAl7mAV8fq6JG86
o4qdw7f0cBcr2JR3g/CVVJHnYzwARYGUCYHIDB9r1maEjfbaHYqdz851TiTu6fLVZxbO3xjMbtiW
7R4LPHMVPZTLrMO+0DZYV3VGh8+uOmfyNlCbWEFM8E+xh+4zylRG/jl1/U4/hSANtUuKuENpS28a
1gOENydUtDQu+JFUU7ZIaJmg/25qThrxMBgck22GL3tdJIyGE2lnDrIQIumF0PMBVxP/Jc/chZR+
hFTqj1K+8Tqim56mIdUahn37Oz3wk1OMTOIJoiHgvthMP7pgrtsiqoAKKNWZi5tGVtd1LyIrtg/G
cr2Zp3q+hyzGuIc9wdKBGUeHyU4Dy9y68n7v+FV3StY3txyB4v+QFzcNWFWjOY5MNgDafozvUAvl
sMnYRLXJJUKlnE0TVyz/LKC0h4HIBHCLQ2YaCNhNLdFTznIsD2zB2NDYOnxfLd5h0Pgd0mH+BmZt
nPaATDDNLqln1Ij6OptSX5gxDb1lAuv5dhKE0RFGMV5JOiY2Uiv2NEA01OvxFpSiMB1w13CBosXo
tyn8QwteaNgN5fTdwc9com/ZI+WqE6qsvCGC+gR9MX4Enhsl3iWEnmCS63QUxdb03AQkQfCDCe5k
IfOA+Uw8P99wh97XDaJp1LhuFnpvbFy3z21db2VY7k4pnB4fzXIJ4FVWaMF8CeN49SJa38zPL7kf
sQV4lot9xvnVgNrjhe1RqgQCjC/Wpk+fjVRVuHYsetTORug7k4t2h3Rb8ZqxBwqHGmizWpoDpmZh
XF+IzH8F8xIslI71RxeY63Sm/QoUj+H85z8VVuv3Qwjc9UjNbz3xuQaYnuKY2k77dxZa0gHLCqcd
AZLVU/+gwdJhmIItPzjK+Fn+lz6FyzndacxND7pJyNzCMg7Yp60wLFiwnqv24vqYCNW7QDG+5FzN
tx2pBsEYtaKI+NL+9Tki07nbl+FdPsbldgy/WA6ji8/OK9t9xXXD/grCUcFVOxaAhd2POfYCI0m1
wQ1YB7//Vk6k7OPCoU6ABIs5FR2GrOI9CU4UrAYbOTP+jNo8zF1FoleouZAVpElf3pOPcDRUhx5I
UoxVShl6chplcU37/tv2vV54rzhSj/dk3oYjWLHcmF0aez2nk5aRGHtrPKn3xgQkJ3dGUrI++V2Q
vcnDDeSut1rru93RWfCsFeddG2BDIarVDFJesJVrPPFTyyTNPraJN9qbejYx/5lQL5UQool8pU9X
odfHVIFEuuo8hlVyzZf1J32K1YAwMskKAcSzO4u1eVkdSPfvM9arTeJWMLHcMPvksQ7gG+hXc3Uj
P2SNzSmPLgJzlC2UI4dpqpgubjN0itT9w/YYU6yFWizAqAWdCxT3kqb7kTmWByqkuw3xx07vpn0B
kiM3wkGm0EE2r8n7xe0UWbrW6D0cR5PxV8C//QXVwsTzZmPpPNSGg6MlFlSxYKG4y3R4bRR0QbIx
o/DIjF4EFgFK/ll4PgdqR7ZztfraEshhDztpzM9fliT6PaIgcbsZ6U8mxatgwkTsZZp1hYnsNo6M
1Yl+lPgDRPE7J/eyFrFRNtTSzB3JrMPlfBjV5YEgzIRzcWOcnCC6E1oOps9o0QAKNT/BtJKwI9PV
ZYBvG+35Vgg3SQ/tlBvM72HQG8JJDCYD7B/IdexizLUW1Pb8bx1Pet5pFF7c/EwlSxoFHKPvp7gf
IWXwxGuuM7/9/EEZjJQzF8i9oRDDdTuP5hirnSZ5qmhL9EF85tO2gtmf7o39utx0wiKGhBfsaVoy
yCg3qF7I7LiyI2IeZ0j8BP3BWVoywOXlsUAEkZpB65V0BicoVd5OGrtDKfX3DexO48Igksednkdc
f2VsAcJN84uWZYIpktMmKuNrUDskLfmgHIQNheft1Z8rzWAZRDdYY3nkiUlQF3SoLKibx2wNUylp
KykDMZlMFytwewvggHfIObOguVmKUSsFr2lYpNou130PkKkJAoSvkKQDnsWTxBzIiHaSeHWHdzWJ
+ebW7v3JrhYV2bRzbOtvv1EN6oe/gLjHw+/pSfmjKBR9T2G8OaTksvFll5rVeK7WUyn1k9QmmQSY
84lo59fFlIIYTBA/0foEMjXkyyhTlKIXJx7JwmO6bjPz2R6R1IaebTX1C9nZykAq3LGC6BNnNFQE
7fP40GcXercztZnHRb7GERH88Yg31YgjlSpxCQOMh+5zlprLpIyP1NiYnTWobQ8mmOF+onZh2pbD
WzBq/108U2q1P+ynCKKFKk9d9ZSE08AZCY57PWCCRx0inLgrDuZ7Cwdse0VC8iTr3vuq5BBw8HwD
7LPgLH4g96jm9I95NO0iF2x/7IUwIDWjL/MD/wty49Rvx58NCsZPyJTCS4MDJtsilgvSkoZIpRtQ
5g4VJO6ZgH1509jSKbuoy3oOnudMmAwdeF805ZzVmSX2+xGqiQE9LLvuOSxxFQIRlcqPW0UCQj+T
TiNkkUh0nlGykqarxUqnOQA7DansWKciH0VrnbwTsExE31ZfOfVglTaSf1GqtgBmYaKKaWVfEVAG
MIt6aVS9gbJBqVwxPlmVkWRq76yYpQu1bH5T9Jo0aOHgvacbJX0FzV20pR9ASXgtnr5IgebVk5YT
08rsMx/vQKnbq1uLNoTJk4hB63n/IhnqWhmZOWOQq88T9IkGt2uLaCXCO7EyDHkN3Ey4Q5bmrOR9
i0Wn8ZKBM72LS9G1XY82f4e1gDwv51JW6eXs6yTFWaRxB+maXLTbKsB5oTsIr/U5D6tjhjRdnj83
UK5T9nrJMuHMNdLFkjgOfNBP4/nIsc76qeTJKkbJDaP2zu4O81VL5nUrJkGcp1PHuSGFJBwXOI0U
/hiwBx9AxFGD9vCP7nF8td/GLc145M4z5NdDk60gCwZ8oW8gDCj+K8dbIbDGhxG3WDbTZ/Gj1xks
DKz1PUkH7CkjkGxK4x5X9nVWsxkMHmx/FiXfXFrEM8co0Y0gZbBr7RZMQqOugn15rhsUGL+3EhaN
E9BTtUp/cp8JmaK+xVToJhDVKlI8h/HN3ysJQ2yXAqw+MM0SUjTy646SMche2zUgFHqNsYDqhix6
vCB7eEHaroSE0jBuzL+fn+fcQx7kRL2IUcXzpfKO3e9DolisvzlOrYdvpiw/44BcGLZAzFrb8a4H
vJhrvy3bdKMCRDAIupwVHpIXzcE75+jvdZp0cj7SvdaRfJ0DlBEl9e4SN7IRSpoI+rjmVkpZm0QJ
HiVUgS/OtPjOev+kf5A2WeBRI++cHL8OgCCI/Y9CkhA4PJajoz0P1ejdQ6S1+nWiuOlLW/Oye3bb
f9e73cQjNlbcIeXR/eL6w5g4YLlLnmkfDD7H08BWEA6v3wlufHok8S+/tVv6nROvf+o/s46oFcIP
Ig9YCV/myUv71oaFVjYNEV0yOJoXc7MwtaO7rBtEXfgl3uhROITI3zhnmUZP3J3AFuyMmGKfXP+g
aM/3Nj3amJw2+bjbuSOkmWeKBz/n+3+QWPo9ioXN5wJDCWA/lU38uReWc9b717QuRC7gErL4sDwn
9p9SdpKMKLC/A9R6hHetngLiURONMmwHlhnjeyarTrn1J+vg+pEe907SFZTtEXZlAqz1uyM62jFG
qqx/g7Zp6QftOA852Etd1vbWMetYb9SA1cXx4d8fWwzwVdhEpGDoJsKZdDtaiJmGRLbXcglx20le
VgnThWhtDaSj0sFlvfbd2SpKGiGOYsPd31A4Mg8rKQSWbagpQ5CZEJWiTfdzpuKXetOE70joI5zP
7wUQyZHz0VCiXNMISzX1O+LWOS9DYW1IuVNHM3rzQ4pWF8Aqe7ZDXeID5krPdsXMZJF3BfRLQGNf
LHjXGqeqMdRPWybseYUtqEhA4tFJ8PaxKsFo97gJLE9Ktw2MnqQRYQ8chnqbuYUBgeYmb1xs3a9U
wU5VzVtFoULhlyJwxK1PCgDQHm6tg81s44OHQRpXEZ07VDTU+B06uIL+jrUFAVE/RaTWFgHRKqrO
CV3DwYAlazL4xDC6lKiogGE6xieJ8FrJYcDlrsTcvV0/O5FQoJbhhL0b1dFDhAtQ7uiqCedNo3ES
Sn8tNGxUFUL5/VobYQL2xEw5Icat2/6EWaQTPotFJ/LRjiRhJucpoYp/FC8AohrluINSqsrV0Rpo
OoSAIL6nYCbLGupPKcYyG/NX5pZLeoT/1CeS3hQxQE/XVfGpuVHI6lqnNNG7k7vpImDR14Yursh0
hLJFH6+SEahiRsm+FCemk4y1Ewi06u5bWj6jbebzhSbkgcMdZATJVe5X9vrBtx1WLpYraPZlc622
vthCOCHvMyCdee1xaO0Fm88TNfzf8IiGQvFCjUquRM0Be8yoJdZPuTq6VFXtAUgFoXubdDMRjpjO
Ua+42X8mtosytnmZ31lKyTRSqtMKebNT8LzegeZ2ElvqqmQ7eBvXalOSox8OXeDlCvd0P5bKcOcL
DhN8pqHuAXdWc+kOx5SIHPLy+lkCwRuo+nGzsuQFBO3IdOhjMECwjejQjnMFp6w4J7P5X3WggLgj
3bppM3euwb5DvRFoVbikJAQu0Iongfu4LBNRX3EUavZIXYbZelcSvIJE65tKG+3Tv0GQPd7svfwr
Sg+yaMW8bvGKWAIIzND8/XQtENoSiJBLY4PQuWGmIJUbgRw841a0YZELgtYr5CdwxYJ2zSefFcnL
d9ARB2aCiLAoP3V9Mw5vaKCf6N73XRLEEyiMWQTHr0rznr/z/5R8Y+hqGvskiUDjA0ZxaX8o0DRX
uj7l0SzrgXCMrS4m79KzfDTuqwdpm3PK7scXhmy/+McoCGb0MKWWSsH2sjT9mQeFET45XCgLJYMv
M1WpszbpAUVbfR9PxzXoBNOZ3ZNNz+yGC+SNOuIxgOhppHFtla/S2gMIAVDPvMIFhHMDsj9d0dDS
HdEajU04a+PbK6jYEQmCBVtQtXNByzKLAHWzZrHr3zUnVgHRZo9VI/4ipxm9zno5F/Q4j4GGRU7q
g56bpOvji1qXZVFghooHLKesFVRmZYIdW4YjTcnHEBwSPxuguW8FKH91YxjdDlxlIjfJmTvY9yOz
RSVAevyNM+OqZItB40HpQFT5K6uGkvH+tBz7s3pKiORdBmKwANR+2rgZafaZEZ7YW9NVjHD4nVoQ
DNSZo/NczlJGxFQ7NgjS/RcAxc8yz5E3gQsxYRiO5oCClmDqn7wSTRVkgrVI3DhqWEHPeKO1mI5Z
kNHZlV8bfjSFNMcANYxj20ufEKjY2Za86pbdG3QfJrHBSCDcB1YUeq94zPmx8QpdPggsn07zTvP8
w+1q6TrVQTQeRW514nYTCTjSEGcbqTUKmOp+pf51Q710bYKHT/pkHOIxGIiW1+4+NRocF5ndMo1c
6iWsf52MKxSxv7So3HnbX1vGeSnq4FPhqxEL4tTy8wXnp4d4zynrh7W2QVsSvI7pudnIu12i+agv
ap0D45XIUo1f+whlhxrYZdToGZ8khWSLJXaTY46+V/k/WhFPYuLzvkk5XQD5iDvsSiSaimzuPlb3
rtvlnIW+0IZy23Q2BjQrIfgoA3CxcM6NHEVjAqzsvOod1zMejz0c6GEa/sfsjc8h467u987M9bPL
BA2dMHY9Qe0h5qR/K1ouUd6QKx9hBMfa3d8r2D4BpiZjm4zjpIzDIacbH2QjIhgHBGjUp0f6wZZD
4AcqHXAhIaRVVcjJxkJMKxeayz6gYIGhdp/2GyqfKxJV5HAGD2OaSfU5Cq5b4uHj+5/JLzIqhTRX
/FuRP7aiH6MLHsVkZKiRX4DzNL0JXsfwd6BuloGbBIxAv19jaYABwwMlg7xRnyxfPXNtI9+UWtvn
U0ERkLbL3PKXrFRlSCCm30aDe9nElXDiFNuvCWPidWAtnzLD2dRyv8hNWRzMXqQiP7rtQDHc/foS
fZ8gImKWQO59Y3fQurJYV7WMQjqtKEX0VYk68tn9hGyIm3VfkJWNqHAga5RKrQqJ5SbMhhxWwsXT
G9jj9dg2QY9gFyJTNWb4PiDoJCiB+Qz25nctt0ZM0tcUxUVtdfAWPrPdApdeBhhPo2q+17W1pMiw
x0b9aUYJxCDQLpsqWQHHlLBYyMAPIlslB6biusA+RI4o2IYveJUKL+UhK7cgLhiFhOWl5jv7otOf
DmPwyyndPwtALQ6qA4Cj7bziFWA+O24FzmqdnnMj1kuaa3nO9CLsNepFDZMKkgXEMhxx+CSsQd7L
WS/jnMl6RGVYZ3sY9gSROaZma40WoNAg/M23deQgJTZZIf0hMv3pvWIdmcjsZIy9dYMoKPyDQpOP
ejpBeioZ9DuJf6tFzdaJVIOCV7qYdxavBVvKQAkh//RGoZrRY9Sa7p8FxAdGRbe4e4pa4mH08WLZ
1TFU8GeDTlcyQwZCsVvOZ8lqmCSCtIoHiC1RP78GHHuS4Q87n3C/EVt/vggC8i9gmWziC90pxP74
+9lWF6Btr6uZ+dUOrtEg/Kpz1CvSS3L853enb6ildWZbxV9dof7EFauXTyzm2VVojjgB78VdPuWu
jJ/+YOWsHV4z5jJJBdv52dtdkmKSJprlrzdikHmv8t79SBRFGq4CXP3vuRdKmgqM4e4e7PaNNWdf
d4GfDcE+JOW6au1maDwf2uGdi42wZwcv/R/1brOupKnieWO5O2vgDiML2iGOVohJtyzeeJasTe/E
ebZYleMOkIgkObup8IAb6iLyzAbbGw4ROongYOMYwnJ23gOjWbN/gT7o0CGhwoX16+CHs+eMjzhi
V8MprhIOd44Ste2BBuGbwZ//3dnSb2eEObKi5SNvZ6VA9sDXQQxjQE/iKHLX95lb13/EcBqweHPe
vQJPG/iUyL5Nu0KX0fWfNFjE/b+hLfv/a8NDjY7Tgine40oTteUidLwpRbVo3J+q0xhmrAMF//ij
ZUG738I9eRZDcEcge82y8kXa5WLwBC6nSjVRIZ7+eB3nCQfz5WAH4PJY7ikTxUCpdmD1CooSHMDa
XjegXEtZOIsBv7Xp6qNwQ1YhcewDw2Su5U84LHZ7KAoqPNFjAddS7tRtxLJBnQ6T0Bo/8nyxa5Vr
C483MKfUXqMhGTzeTYbgqG+tjYVRTq59ZQbx2KbiRRPmF2WmrNpVKl4VyO3+WeTKK9/PcIY+Lmlr
VdWwA1kro43MhnxZsDMeYUUXrEFTLywHt9spmPKEKanTnVeophs0sZSAqJkRb0fdq2iW+s4H2W/A
CyFbm2WcM9oz+8uMqGiFW2D8E8nFYHqJXr5hhG03t25vNNjMJ8j5puBnPcjZE5oZyH3wGkxVggRi
hQyMMRFRTUhXBdGeXJr2797q4W09RdfNvYlztLPXBMwSDeKTTUxoFhcKMI2BJK0F0lfaa3wjU15j
95cgtp4Q32OL+5+xYtN1ggOFQS3X93nYQyzdr4StGRdVWSt3vrNcHjfI2jW1HUp4hB9Pa4Sz0L0O
//wnENC82EUZedpi4t84GapPsByjjD9mQmVtnf5aL6TLC157V8K1uJPgRvl3uJykavaxuMHv7pHW
rQQjo3PRYq9PsIGLuy49HakOQjZqLahsAmi440EiypVLoHRCkCCQ/dNppRmB22E0p0ePlRnc/QC1
Tu7lbrBTug49gWf8lNQlQQIKU42NI2m8Q5lZXphWdmGF9uXQa6ydsCY+b5MlSPCtHPtv03FsabXy
vlVxqFEig6RRZ0JqdUK9yAAEiP/h5vT109YPdMcM+5ki8Vwqfcwr0j3x2QnlQM+hlLGDXqP8Ayl8
P4pnyjuuNRrL2cI0+2Y/LNmG6iWTaUR1FPnUzjvcgkokE+L1OUY/Tw+SHEFjUaBCLA7hDp9L2kCI
2Mv1ZjY4APCMV5HNMlhNBtI+nrviZr4IEAhoYTE1XWHDxKIaKZx/fNJoVDRgiNAIVtbNTRyRGxXg
tR0XtuEGNXTn7VCqJFebAv0AFUIJ+NWto60fkzebHzB6j+7B1vdriVqNln3bUL2C498gUNDCjRqq
4VycSHwYZhURiFdq2J3KmJ5QSDoM2PB0E+hjEPnfeuVDbOE3JayUgc/4ZY/xelZOT87VgHRk7GjT
hdHotK/ZRaDVeRmEHBCDCB7HH1uJMIv91F0TvWiImSL4P301yf/avs/3CMbjyElXURgAj55Uklsq
3WQBGTKWzzf7/IVjMxT5eyAd2shvqezE083ck6Ly2AET/cCXLnxboAZ5z8NC8+2CJS/LzUxtCUWS
MY2j75p+F08BOWROUXCoDYbueF4QPvp5GKRiaoTP65xV1Cn5es/PWcevcOG0jphDWQms0vP0CfDq
okaxaFDKo7LIWtA6DUljf7METtRGBcGniufbRq2TYNjDmo2PjNDstA3cGHtQavb4Bgv7mndT9Xdx
Mf9WmKHeW6HrtTpbUOnmHnhgO9XBBirFjd1fDw96LFQAUkfFsRm0QJ36BSK0FTmQL2Rl4R/FL5TD
fkN9UyAukwH3iGjX4Rkvn+dFF7KAhdEl1sEsp7TCy3hBJp/eIUOY2gn/ha3o3dOLL0vS+C3N+hWK
9Gq5pmAylkY2hEW3sICYeO9aC3t+93mU7Csm0fnLP0dUapLIlmZ9OR4soLIN8ub45E+0Ywe+TbLY
noJmKB6ygxpqUSMm6aL1mLVRFN8t9S7zyUAqj0TQZvDEio/kFDF3GaZS+ePXoVxwTsqCSJ4zoGdm
Qt7pmI71YOv1s/+8WLuoZBkREUvQwUMARyno3Ityj3g7GDhKpXc1B/9xaJqZ1yLch23Ek3mMETXA
O6DULCh2EA71q5X0+qxgk2nSe4daDe259POigEyQDOdxYiw0HZCBG85z/sGAh92bvIXfRK4JRUiS
Wx48Ur8C9ypDxoVKwLYbt4g1ZQiwq4J9LJXI/oXPggE+KT6C+e9Uwc9EA17BgsdeWe0ZeqLMPwfl
S8G5iC/GfyKGnZpJ43QP5z83G0z5cQFnAoIobvTtSz5jDo2+x56yXeb09ykk7MGSfz2PTEbOH1pX
XifEP6oe44Gbd/HjAzF5L1XFW+rlw4bp81uS2Lm0Euwycl+3wZApy6FaDbB9uxF2B1q2zQEVBSXo
Y1l/uZfykaPBM37ltzOmmS3fWrSARkEcn18xSYuRJLBJyk8SeRH8T6VQQQIOfQn0XQnIx4ANDd7i
MsYSoVSVI/RocjeGr18C6cm+beejM3LWGipSNhGfYS83oSmqKxrleOrhWJRFXn1wfBZikYlrslUq
Uz7BfdXkCp7C1EZbQYYDh+lH4KCF9sjmLXRguj1N/lgSv11HL6tmIIa3QyR+jJOTjLJqDAna6+m1
xYtAYvFUtnnHHSPsbLS8DOXDsGWeo+DteD8ZO3yOpAYbI3uVUO2bzfYIX1+wZj8iiYoqX3eY1tmz
MC2FaIE5iODisUQqFJCH8r65Zl5MEglV8QMrog/CsznzSG99ha+u1vy5CfavCFe5GxlHUuQEU0dJ
vIT0t+O6YkSjZF4GP9CrAp3rnXAXIKrxP+amIppXNMdzPuywOugdLUNZBNbc2FBwLTu7rhESk3q2
9leWzaui4rJdGWTRkm9h/3J4T8eg8dv1z6738eBJyRdI+0IO5d8kwYbAB8JnS2YdHaeIB/orN4sZ
dMTga+DuwZn8fIO5taxgAUyUfrfAUPG9vfGDgysK8I+iXvVpjivugm4GQD5zLG1jEc6TmPxTCZ8k
y99qf1Z/uwJrTQYMQfMtq/AAB0ZFWO0KMSZUeIvBnkP9TgJqmDJueb0LRxfX0O2e2tWLc8pFcoTF
NWBESYuGJpOvniKGX6aj5MdxPS7GM6QN2kQlCzPMHPBzhAV5Ph7vx9JG0/ZwZcWztb9iUs0ox/+K
qG3STGtKneuLaDLxVqclKMIFgNNkvq7kn5JdkCxxIxc9e+RjRAy2ofNl6eMFh3/tOX4UwkXfb2JD
EBTVts8kQd4/HzGh8tOdno4Rwbc7HmmDK4BGx/rJuUBUsNGU392y3ZydGnHGN2FZ22iaKwvMhcnP
hFo/GYtlG6Pr7KuVdVM1dXfisaf1r5TxvYB8L5pjsJEMnGtZgCXWsL4Tt6zQz5Ji49n+5SOMwfJC
Y6sQ2Muf7MXPhls6LTap+Sd67/UzLKSmgN6UzswbAFRAgGttxDMXlfWamnymTOHW8dxsWUYSyyAD
bZ6JUbFx//wG+SlUY6uIhhmQ0Kv99w36U3X6BGYuI4FPe5nTKqDlB7UOg5Bguv1jvKEjR+gcEMmO
+8JMtNPfN5GKiVF7xhEJCUNHQN/hKtbhXHxtnGmAFmkdx2ltR0S2EKDeEF5J8+kS7UeegD3m4p58
KgFgxVTWWeacjvDMIfmlcZdSiEh5+NLxIRygCAKH83s3UOH4jh+QZGCnfN7RB6u0kNUudB3VOG6V
TF4JnSvjTKUNeSWCjOYAjKzVkin7nl22KEZjijRk+8LhLChriIYVeqUExn+FP0uZhuJVUS5jXf37
7xpQZ9/LT2gqoLBm9jBsLN11WbVoSnVsYYEr2XUWCFmN8NSJV/RLiOj8FgBSDtUk2AdJrYk/N1EW
jKVoWmTmzPsHO4zzTebf1els4+87F1+csMA0YtRJ4SLkdA2OoQX56JprvQ/4fxQaxZp9/FA9jNI2
Db9A5H4hIYkc/PGyqUS9NfNQjLRXUbgyOWwBDjTgxMgnHanVrVZce+FUiV1icvsYKJcu9EkZz72/
vPOIP3P1KbGGlRi6G6xS9C0pidcDRW3DWqbmCA87TmjGf0MsqEaDG6fg6s+WVZvQrQLdhnqT0Ext
nUKXpUBLkjC0b09RqCmD1NXxn3lT+Hcd1CpzYfzNOp9x1bL6qNKAoVy31gRDGofMCQMZF4V1ELza
4iQss3+dy462TIZM7BmozDlgyX2QydM7gBClmTIOH2leXkcQTh1VJOnoSyF1Ab0jE8xx2ImTOjQo
ygiD3jBw9y2K8EHHpLm69q5KaQvB9bf+PnwXko8+eoze5MoPtyYFGKKjN1RYbjtqINL9IyxWRWss
PxocX8YPcAwq/cRg2W6Yh5WL5jBAg02pkIbf+gV0ergcRmRr1ifTl8Ht9N6NQU+xADfBaGo/5nj4
5uNJVKkRRC3oeQkufhpZGNCntpeqYwQgpHFEojG3Tm+X061llL28QVGfLdvNiiXkG82Hxv0O8+No
jgXLA08dwegofi9s77iVHC7cc98ZBznsk82XdjvUDkUZshzjsZcApfJzQBXTo7ahsTD3xVkAnPtu
keP2sXQaNWh2tJc/yS0iTUHdK39wc+yV1f3wIn/5TdtH3+Doey0mbjMxpL+DI/Ity/C2q1QuX7NW
awKI7F66BpVoPFXTas7JIXiZ8siFFF1XeYhjSz4n5NTr/JFxIddZX2tWI4aAyojJpw2/VqTLb/Ak
qSYXdapguYqEqN2qamIty082/qWCq6sXl9hTQB0s9MJBZuJ2foV2SA79lM1caxos501fvox7/zWk
Nzve+KSoTfjfkuVUQ1QlKtmRKX5qm1uOMVwCCNae06ExpYhgL1vvNFmQf8mfGodygH4UlGNfdweI
zDEXRF7aSDDy5g+kLj6zaESFH+pdmz68qa8ryNK3q49+QXIP6QIUsxhf2hGXmbl2XrxtUgJsUhIJ
2Ux+mi5pXr1ffG0CqScAz7sz0CNUrhOGmPKpEYUY39vCwtDE/dzMmyCDdqBwQnsmasXnCDk/Onlo
SWL2sYY2L9Obiz8lQ/1EER8rGMQPjrKJ6gZZ2OXG33JLQ//VcY28Mxnmn+0GG+PJbazEZwe51aLU
DAxJNa1+cpwVOYWHcNvJ2d+/DyhE/UZAHjtXzZSG7aTYe2Q9yeiJ4lWZt0UxECbTMcBL+ToE1+1c
hHmdQNCrsNj7kFfA5qxEz5PCxK5R+eSS+KAZAkfDKxLSTTNLenQL8xjhE0hfb9FD9UmcB7D17ywK
OVCM+3awPtcBPVOZTTMuVlV6cqxmChXqoZSFeBOPMqdF4olp9Xmr1ZqO8gOyQeoYFYbE7y1bSt7t
tJNAvIid5vk19400ExwOJ1Ef5cqPv7wuLQfD22z5hYg4C6+RZrep/GSKNZhGwHlgTWBpwZvssLUf
AoqChtKuKaj06XIvKmo6LLzifQUYxMLlcS/OneC9ozPS5VUVoafvxzNbBUod9og4A8+5ovXPSAlv
h1taEh2yMcpGESo+yOVQofOKtRMrL4Su4bMUt8PxBhWprXokX/EKbqpLmXitLmYvyF3pWr4R6KPV
1R1e+ThKjhEJwccNkmO03TlTshx4mD+jF0VoMc1ZvlIztLGqOirDV7gg5PU0BgJXyDIaddwCiWvV
wiIfLDLFEh9Yib4x1fVeaiw1fOIv6hPoWdytSg9HumTaNF0xAloCq2ik6k8qukphdI8QAP4wcdoE
XEKjYHvM95LZT+8FjGkj55p3BKut3+iA1RPA4jCPppPEXGO6PzCEbM6uBM1/6Xd4esaSuVrYyRHY
u36aLRePkjAamBw+FhlJKAeiD1kqhK6fnXbXxYTBSwrVGcC3HJZN5f2QF4BZE3FphXVjTqkNZ+yP
iRph1g/wddZS1a/mUz6tJPeef9WkJ2PIfpqzQIZlCpzVcafzL4VnEbnif2tqMJzaTLO69CvvrYrN
r0AigR7ETzsANUXlCwfhBWeQhTFuYD1ASaoL451373n4IikV4o9r1g0hxdZAJP4JZAjQ0eNtMwtY
iD9RMoPX0xZ14Fy9zDWrx4HgrR5Kwe/Skj1DrIhE6fGdymeMqU7zqMMuVjHOAeGMpSwSgUSehyNW
72y/kWqQzbUJXJXG8+q54M2YzQv1aP7cbAaQpDMrqQNOwCqEPs72J5XHJXHD4k2SQa4Ir2oZF2Zy
+i58ioC9AiaJLFLZtaEuzyZOVtKAD9emdtdfA2rB8Ps/05hR+7LyqZlAsPDzE8ZszGUqwNC+oC7W
xCk8YlRjMXvlVn0RsWcOE6uuz/mxYdv54fUYRx5WeunZcMG+2ed5oFLHb2lULYwboj77xP3+SFG6
1NjO3pzVZxHop/TCOH5ChBd8Wy1cy7drugMldebqRzhqmLjJo5hT3b0WLpLq9QFxig/c+TNXuvzl
hBaZAymwOda+uQI69IdPCM5y8ca7PaE0/SNRiztBQ+b8bAPzckrj0nNFGaKXdEGZFkUc/i4CkzAx
hvYFOjy9tiCcBWwcbe7lIFnPeJkSZvuF4XSAbl8eqffCEqFoHjTEEEnn85Nm8/LSdWEv3xezLl+7
ubtlGID8Yp09Jaa69PjH8VTYACxgJdI+YtzH4G1hXTT/ZtRS4ddv8EdLhAf5PthBYsVYZ/DK4v+P
+cwc3gLCxyC575HNHfueVjPV/TjvU2CagF8pobYJsQdPEkbwmtgR5nrJV6x7hc/ntyo9RyQgzlPe
M0Ngmryq510e3eZe8vzln3JRAdvcJ947EYYrxPWrvn/Cyd4Ia+rq4W5XRgSAck5HT4ZvfzMhlMJp
19iT+gElkQxYyYZnJYvGM3Et6tU4jOyYUFFT4ROuRT4DVmSTQI0yfnuEQv6G8tbsT8RBE6zWTrtP
3sYrJUg2024073rno1RCQ0vh5dlqZIcRxIeR6Y7jCJN5/yldOJBBuEb8kwfsD3vhEi0qXd5zcmoU
dPqMUved2LlPhfNdb/EgErAqIAb2KPmoeTFuT3jZzWP2uePpvQgkPbd8mcJVlGp+uO/nGE5ECHrF
MXVZS/qEhpM03SsRwErcxlvbfIo2THSSGM8Jr8V5ASm0E2O3JpqR+17Hwip6DKsfq+2MH3fI4j7c
4ZzLQr+1Wi2+jJpf1k7IBa583eAviN3d6F9XdzR/jY/I+7l6J5euca9omJxzjlJ0uJXukdJYzh2p
Sv0yruEC/PlkfeqcS3IsHWND8xhykyHvFFgKdwMpNSeL+u+lcsY2nzGBs7q///vbs54cCEC41L08
cfSMzl1CId+WlIh7B0zNBhbb7+U+yf0JF9BJsKp+4t9PsHivbL8FyOVQmxlSa/xZPNCfCX+HZbeK
xX02bRYkFmDpiORqtrg11IRuzYo2dgf3cbjzGsFnSCIcBP4mBV/WxeZtk6m+NfcLhbrk2881gNZo
ieaBTXpctjfuBNBscKlxR/SC6DbEceWF8TAxi+3vRIMxNjwOf4lw7alipesB7QCRHZ26oS5eEIhr
DRp7MiigEZ7pMtpVIrHT3e2sW7Pd5MJUuAf+fQaIPxzZbBg0EagEWwXoREzIVwMQxmGfPnZAoIdm
mp5rSK853B2I7IaGbBqGQvHJyDUn5a7B8aggCOdQtQ2kG6bgh9U28dpq9EdRTVQT857iJ4GdqUsn
cTA3nfWiZC3IKbT9WiIq0qiryBm3NwWP8VGYUY+XV+8LCSO3zfeUEs0Il5lFgcSCJb6tSiw7RHIR
vxiTXOs5PLY9NDc7r2JqJAvJ2cJzEv2VoCMJhpPmBvd0CL9aEQtNShpqC4mI7VvyV+DShhCKd/PX
XLbQca+ecvAMskCl1lNl+lmSrnZr8HBxCcaTEu3fm7sSlPEndhRUh8obRf345ULim/+Ka5dU2AWA
gIhPVu5bueu7BKPHFLfusRSOdCDfqSW7TNue9cwC15AwoR9S9CnyQHi0uwQQ2yzPAkZFTvO9xIc0
v2GYbPHsAxd5pLKDYm+B5hzLDDhrDNaSQBK/pJjEYFNJxlEFxvZjJqaETTcxHo8deDzQbcS+V3xk
gipFcE7bNwa1U4L70J+N5xIkWL/jLfMAyUZ3o8IkV47Dj5NliZEdLkyq26CdOXC1PbdHAjPt0P4d
+DxiLxGAFOML6deTx8xN3F3LsdsJM0KMVY7jvjIVOm5qIvNyvzPdZY874weC5d6YuarzdHeVrt/Q
6kDdOLDkH02+fnY3SkYIe/r8XPoiIpXnkBJ+rFU+raFg1ZJJ172Ixqm52pF4RRCAcobQiVBbaJj+
6Ni8rtptmTZquuoMGTkpJehf1bne+UE3yKlBQeFC8ZrjiDstZW1BDHcTaepNWFUs8QQY7/pvtF5k
mGW75pZLnc7HRmvdh1VcS+Ne+YZRVaRGDOjqhZSljhE7fixrYDkpb8PY4Fn7HIc1Xa06cgcb98ja
np8g87RULMgiYuZ10xa+/yhXmWovBi1o3bjz0A8Sick4apAH8tToYwbXJV7dwbrIfhRsatGEn6We
arSnJ0iZh0Oypx98X+dIwjsSYcpM/QRa3X6rsD15P412/voxfDjivxXCuMf8zvh8VG0hMmBax3YN
zyPo10MGazryBcsGXcqW1cg11CDM3T5f5UUowzOcbPToBErUeFJv47xvC/BvSgTn56c04hyS5wOg
ttdlqATtXASMuu0o3ekaixsoESlKXie49iZB3juFKm7XtawMFyQjHZnLsXp9/lF8a2jUYTVn3/jE
fAVKI0EW2qJN7ArI6OiachFWE02HiC7FtqccSsMnW93Y1juSKUXT4H42iAFNGvCSLHhQGNCsQARA
J9mDKRGKdTTMkb00ob5tf5nCus03VHikl71b0ntnxOY97lQD9jKNmq1w5nXr95ckKuDm/s+y9GG0
txr7jWzmIT5aSqEFzgK4MoGadBBl7j2gGcVg6q7V6eKWRj8asPylJT1rboYEWoBmkCVoynjyz58A
WmyNuaK0fGwB9uq6hb0ObODXbXBjwjfig9Vv+ypyKXLAe9XYsK0m3s8PU0aBvN0EP/lpjNXDPQaF
oWt71oztZ1msrxTV4WZHeCL4Fv/RZD/l6des0dROT2fxlihTBbsTvFBCVMGWg2TlaEhqlO3KlgwW
8mlo8fWpONUQg9Ax+qx/nXnLfM8pe4LEY0gxS2dxOy9jjAHM9JXC0swYCG+HB4rF7Uv0nnzRNyUi
eV1YeqNzI0VFz79GvAPwnM0vGAWAwnZ3RYAzv0OGetvyxlKPr4H0cnw3dyRMnzwGYBqKbygLzeFl
K+kPv4qbkItZU2Ce5230p1ykXDEULuVJln8U86gMuTxF4/vMQVZMJ81osmE53Q74lBEdmntuUrdM
Ba0/+scQGhEvVrRscG7TgeScqvWtsR5P/tqVdPiDcv6uljR3Buhhg6MCwazKz6+uw3tSIA2A5NUB
MG5Csnn1zuO/hzZtQCzFvQ0HjyAnRxPymBiiaurMiToFlZBxYysgsiEfkLZjPMBwiWCA9CNj0TqU
wVPo11e8zoy5JPANLB72dqKyuH8xWpLPeYFhcaiB5i4xIgqkT58+FoK5at1FEePmp4dzDjx/UVTl
g+XRlMhsyYqwOcMQ6vxx+GjWh0tcMQsDMiKqBqJjBFq8oF0lH7SMC+jfsoKecOP9AO3JeSQuaDyd
edeonFw4TqgyCcIByqLADsXiGej7ImJ7Jf+hnwLOdARB+7TrAyVJbwZxrHJ+jkhDcxyaexelBpB8
0qKcqsuAJZPfMQbE+ahNwWi4iB6sLHI/WFMYObWb+E3FU7t8c768FG1z1ffK1uGavkcS0+d92noS
GShvD1uDfnRY0ubcYpO4WYmJ0pdXhQ3mFnGMp1oYfT2Xdew+CfqATMZ5RuqYEn1XJTmbzOxX97Rd
cMfvwzO2F+UuNvlWdihqkFCvbCTNbLqgjKs+oXdURLK2OuBpacib+2zKenrWeR1GWJi+sNiLEQWM
V7tVefRHYxh8X34aaijCK0zvQvj7+EtG5NY6J2V1TduedsWiiTuXZbiDy/gwzkiQjhxF3TFWdyaR
U075f2ujolWoVSku8QPBI+IF8aVwhLJHRoomjr4RFKgs3LAIdvywdwNvBmNmvmqUzi4fTFFWDFUs
p00nM+qwD0ZBuDKfFADcNACKfqRmpsV5USdQGaOimqtMe+HX/hhQnvEVWOQw1MVNYdTG6ipvu4FW
lm9Q0hKXaxq8JsByybWyApRBOv3cKCgGD4rn5B00q1IhEzGCSaNHj0fFl6He6silLoDZo5SCfYU5
uewwb4eb+BHAVHS8brOyMc+JhZcJ51OFJu+urgoqxz91D39WA7QOnO2IDhNkx6SvehFhxrFBCaAW
GcGmjOBNopkYxn3pAt60Gb3qIm6Eo9NHEWLrI1VmPywqjzNpT5N07cJ1jmq+zy2DXg/9rg2vCsXK
g4FCYil1uvdyMh29CVmCicvLUkZ51Uh17ybgOiivi4fyDrRXLgkmRCr/jUnVwRGr9dWvvK54gnBN
sWJ1oFlG/NcWcM17cYrXpzwrlZEWMaP11EozJGwfu/i27+AM45h4Nm7jeiUvRmRh1gzwVtP9XtNr
afNx9THuQDBk7hSsN81cAM75RRvo9P5xQp9DFFJy+d3ydE6b4mssTUxJOH+MfC/cyJDdE+MbLYPk
BlnoDiguLRQ9HhtHx4wHfC+BNhaqycxPsjBpQOkFRru530woX67PwfxLT1d2EONzxkig4pOn8ycL
K7CfRZINrd3vCk4sjIFlygqGV1J7M5mWwJ+FebC8BvgO2sVpHZQ+Wk+QOIxjBoONmfochmEk18l7
bFvnRMjsqQPS5dSvcQNAyH/qIBykmBxfnLlnmkBDEbUBg3iuexs3wCtEN+yEcx27zsvdAAC/px4O
TobSggYoxV+n4L5GnS9dRN2JbixhZM/1NP0y+kD9fobvxgIpu2Y2OmGBPiz0olUpylRgfFjyUAZk
W72CTC5Ysa3HYPkyv2zMHxHp6YkIYWVotyfdK1B3aAqKWyw7SVZ8APkFkU+S01C19CmE6UHAcduh
edHx6YrFXeF5JTqJGmY50bS0zZqTMMYpSYDchBLcYyAsl2XdBE9IhmD0qjd1IkkqmzK7iQwuEqNi
H/nJmplfcadjkChhZ0HxnsSCLrSiQDkGm2V+j55LdSBEF89y8JxPwsKhyXubxHQ9do4Sa3oJFxyv
4O9+WPipDSzJ2r92SY1mt5/zyNgSUAHvpBLdl+Nb0W9v+5MaeNdTPqiYUeb6f1gErJmwzMRzrIBV
/G7GdZQMd779S0vYMQw+K+klFKPmEQwooEyy4tZPirsqiVQqRy8rF7i6PRJd35wu7hZbWyj9ZXbN
d6GJHLjYoJKQ+zkXSRklEEgVOsLJkmy1eb8VUbcnalsmR+t6YBcwNFqlRT2y0KC3lPJcnL52cNP4
dXs9JdXQNlGkCDdzPcdgs/3+BaPUgyx9wSwRhX3JQVLRgMLFr3ZlUgraaQOerrGHCuLY9JLtBX2s
y37Tw2pShbDZj2O9FMcgzZ1ENV8JIlG+lc3R0OxRfLqAdCiJoOCxsR+fMuCGdHb2cWoOErwO51rn
r97pTDgZhshLczYPHRkucUI6az2eyKmoNPbDn8gPJtFlBYqVc0IbN+HMswo3hszhSaNc4KWhD3hN
gwHNhHorBMsDG0yHbykqJFrlodQCuLTfs0FyN7NnuxpKyTky9vPP5DxoaIr7y9kJpNgbKmYyFxCl
rG1sYphH3LX3yQ7bLEdwyEOMr9n+tadUWevjTP3YuQ+KmEV6HPiyQnDBO6oua+aFj6ETjW08zVMZ
ryhxsCJ2iKY1WWYVk9GXmrEli/VSPElZeymSQdsrTT/R7SqFBXqhEgWK90t97PN7ODoke93aCVMJ
wdSrKDInUAdVb/hfnxVuPn1YP4lBS41m04+gCNNrw4rs5DGDrC10uKge8SXB/0GiwztUCrmBONdF
RE4e+4pAI0kQgvtzCxcHBOvSlEkqsFNVPzpCrg818MCA1vH8GKYx1zPzIheNP3vFFuK/pSPZ1oRR
B6a2J31r1l9YS9zYH2hTmikNFypywfUx3YLeNmYtf6fJI86f8HQ/ADzUciyItBd8EBesD9KbQuXR
1GQeb0gYI/SrEFFhz2ujD6YGPNqre1asXXjquflZYrqWA7bm7dtSsW5E3VOtKPNecu97Buam1pRE
3Cj4gnCz0+7o4+hdAbS8JPXfvH+xY3pwV2JnKUl/6/2+C14574hnaxbPNUkbn4LPLF00DCnu6Ovq
azRWOt+zbPauvTOihxxH/+fhvu3Br9kcoADN+w6Ia3RwcEg8T4vbmhlo/fjhnqHatxN4S6FxvKin
oiCL1V4JtgYo6iO0scDL6v0mU6zra2aVX748rKLVFndxZmaFOzE//WHUeNzmbKZ3O9hr7Muz2Fm/
ar2y+kQG39lv4dU2YEIInhRYj93I9R4RR9v1n+pZiWUvBL604oXY3UZfgC0GTtSNPWz9kSPzWEjx
2JnsstZBUA3hid7CsR8qJrdsvp7Pk1wvcOUNPe9l3CnXxIePb12rU4e3WmqNPLLZI2HX8CTAPAIw
5hbvmq2tKKtNjx6+8vwnhA+41IkjBwnY5MaC9yLXgdyLr3bj9R0igjYoAykYY1CigcfAwp99q1l1
vIYA5qr9389o3PBerKWriTUpcrHdYQQjInUoUA56WK1AxoGImqlq0kdw4l/z3/6U83sY9iMJXTeJ
kQI1j2Psc0HnObO+SGPJuvm8w+uKeNkAuz3Fbf9KMpAtRtGEK/QGJitJVSDEJ2yz1uAeXWyCrBpp
NM7J/cdlDdHO2S/UgL3DcaxDMDnMzU+AO0HSRm2d8gvUZu7bYm2Z7JXNeHI7SycA1SbftmgFv7NQ
sVygD+YwF7nsLIug3FsWHHfrRNmWcw0xb5fyjlkkzEdf5qTJSj22Ol+lRqL98EEjWR4+8aP3PYCs
t+K4zAhm3kQvjuOsE7rZvmrqp2mrD5FQuAchDGr3nQYzGFG6/68/ne0E8gUrGzZSs1NcDPXjPTA7
lxSNumyi0LJbxpWh0fwFoTqT7MDlJwlXmrF9uEYNPg7MaB6l/xjf0QHL3nsM4+DHU7QRlbhRq40f
Lzx8+P1h3INwfUthom6vpJgUt+7NfUCBOGh9b7DTxrIE2TSVPWEaaNiQVhVgxfJ3sF5eSMwFZS1w
0VbspRuMpeOHY+PJSMQst3JSpBJNHo4Pyv0Aky52MxfG6mp1i/xOrHiTxNhssOaU2D+++t3HxSYV
fCfUDA6YlYTvvt4Ae0K0Ri+H1K77RklyFUgom+k49rp3VEqRdtvHhqsojGbqFTVE755BqXfH+49W
HcPgHjWn2ocCZbj/fBqP+vQXUnIQ0pbL7Jt+lIbxvZt2a8Ocn0bz1XiE2qnVlZP0pbmrnTn/xJ4/
1wCLjMY5cLWznxWUzj/rVNbaMN/xPcNdQpb8Ow5C/iA7tV96XfW9ejqh0I9SlL07Dl8At+xHuNR4
97s4HEmZB+FKuDyYqCH20zMg4Q7UtSPCqE6gJBDotdfh51H3SqkEehqFJSepp9/NnwhRTE2phDqU
KiS6xXgAd7gjbK1pdfuogXBKte5gdPF/whhf/NQw2ErPMJ8RnE5eyIacKbt4OE4/6Lk/F8MPjDwI
kFfDtHyL2YBJH0NHFIB+3gRd4BUnKldT7Qn2OvWo8TdTaJBuF8dJlLkPC3efNr6VPqlWzIIVfuRp
XWL/2+8A2NCRhFNjZj30XqmqEWtpNec77jWdB07oUYrZbqrowvlAot+pgQrD+F1LEeSBmPCPSlEf
lreiqavgCoZYN1hHyzbkkDA6pUD0IRwPc3DVMFXp1OXeqSd8UwtrH1VNMdMTzQ0+lvYn/ZDibUa4
s3SanhviWrMLrO0FHTNYmekljCqTouNpZSg4eTAYKAG6FETxc4tkfgcY+zhbhHu08Q/3z8lCVH12
p/e52XM+mNNixvcPdnflqxmy+fx+QPiX7s4+NyHattLRNw0SwluFD5PHREQ1X1J17AbOHczpQDKy
tC+Jk2vzpnCvuTgo4euB1bR1hVvQCNkxxsNJ7pJ4KTP+NcS3+OCVH9CgOsLoCViigfWU3dToVMP2
NljC6u/9anIBV9aikAF9Ke+VRtT3unL+yZZe5xE8QQ0T+Ll0pi7mNfRvCi4wfC0fJfINaoOvLfGX
7AaD8ZoVdvy2LB7nN8Ee51UU5Xb4yYcDbEDeGX9CYsbJ1R3NWFa4dvpQM14Pe7/2UI9jVGTneP6Y
EjZPi8JKKr2DWTJFz8p4+UliQrroEcU/Db7+TVdKW3TDxbfLDI8aTElU3/RBQGBwhKzQCzRH15y1
GYQK5yr3WKbC7YNVaJg4efftehRReetnC0BRpM1eyUCMdFYSHx8DKtjEbZMR39OeOvMGae39k4Ww
V9uIMBMD2VEidNZf381L56fd6E1rBm6ke94I5Ptpo2gwCF+pXU5flc1QlugogvzVF9Y9kZT6N1RS
EGXKIWQiA+iGDons9QhCofZXmWbVMlbuJE8xzNhGON+QabVJGPODyRktn4jXRmagrTrP5kAWGv7+
OuneJYXhMdVefsZ/6jLMnfyR5EqLD0kDIYxejVxajyj7ACpaOFQi7nfv6CSL73/6rk3clI2ZCEoj
WInxRt28iD+Bui17/aj8vdf5VkLTiTicoN4J6YFDJltIUOwsPnZJvc74O3hD0Jq0VGJn0mo06vCZ
/g4/Xgk5QuG3ZXkNxnlqZfIdWKgZhM5AiUWsq2qhUp1I6//UCZP4NXt9+U71LnricfUnA1dblGlg
/IBMhSPmNTZdTp81j/kcclmnO/62K9YkguIxr3nb2lRGWrs+uo6OMf6om/8pB998Z7OG9gN/MZg4
Pvi1mb5yALSCsiFkS1Qn6uG4lyFxuxHsyUPPAIpbiHniVOyt3vZeDhyM1HVTfjN8K0v5At02JOKi
v/i80kt+9khIj6RQ1efWxDUmiJdUqb8EeyVt45Da5FTir3iIoN9iVexm26vuKlG28lHvCQhRWETY
iYsws7ah6aGMGpu7T97VivtYtJ9VzqLnE8xPjT2rPC+NlWSzEl5euoCW3CjKN0o6aAh4I8uti4DY
kyMZnUxq8WFOfXvc2rEm70azPvrxHtHaL7T8UXQgA5PIAeWPktj75FJjlGHInaGIadvBjkrQ1yWk
fIH8NT0maY+ZQsgJDvk4RLKEoOrO0vXGtFIfNcMRQQXnyBp7SA0szDzgzxJVqSYtYASX/G5OR5Qg
pnr2AbB4mm/DiDd0mhDVBVx10Q0kRycT6iH2Wd239fz+vO8HjnIR20PFJEB5sOU15V9VuTInPcJc
8bKFIy9IeCOIh2HZPO7nl01UTKSuO8kV9u4ulq+UCNtAqn0VxyV6v1OvaubVnqvAfKAn/g5pIzEx
LR5uLwP2sPTv0jFzut7t3lJ7rPaRomYKbNv1nPlO48e4wMVer6u1yQk0UdCY20QHVDJ+ylksrem3
nsFR6DPThLkrXJFzLMdt0BOiXGVZEDeD0KQOXbPoG7KLU5LmZpOKCocKelCKA+nNO0Vx7O2xnfw/
UWAtQy1xyGz923QxccklDuIK878Zqb2OqgznJU8ncs1rg8+zNH7GHrYEkPFUwyXeIt7FXAGFoXjZ
4lnkk9/sBfQd2rlcioy5cjwrH7rpWlBzI1Adrk3GaJAof1tNu8AUMZhMVpFIYIJj8QAXjIQ2oNqa
ZYKx4uuqTsUSE0AjEVvV7FXZYR5E+Hkrfx57USERfOR6EVpIOARBUY5duInD59LDMUSnOWawTgca
VWHc5jtRulUdnlTDeWkVZ/dxHCD3A+Z3yBGcsUK5IVmu3UB5HEf4c2RaOeYD5wRUTT/kfi5/GyZ9
YD5t1pDxxWDSRWaX3yeFJcNhcoCHUpDYOoltS9hcAj9u1cgTCzK497ErKf1426dGlGsQ2c8daXyW
QTuYurklmxjJHvQIzmJPXvZ3/w3RBAurIV2NAAz0x5xaEm/F2dJvO37wnzeq0FIehyd80bzDoV9F
bDOkuuh+1OV+eCLUU48Lm6MInE6TP0LuhZrKWh74iImHA+/2Dz/CGHYQXhY6V0PH2lUYTjwJ8OKu
069n5kJM52oNNQL48RtfYHNgN4+wMdfvVmOqTDHAh8VupUpgYsskWqS4nJXZoT/FjuF3fYohvMSV
Ag//rXAy1CGo/DQEM9pHw9AlqdhGqnB+Y+dW/ppU6VuSWJkiPUiHSnoIrnuTsbcrrl3qlHt5LC6/
WFe2Qi4N3B/OGq7icxpCrB44YMyAIsduj+Ly28yoSlIVFyfIH30BdnZgWocfVYRixSS/r7AgKYma
srEZW35Y+4FK0QkopQV7OOnjmiBADQDPsIvE4fABYI+JJBACWPUh8OPrj0xxclEvtWERxImCIA3K
g9c47OvQg55Bi/Y1AE0C+C2/l3x8tEYl8EmXiLknnE4POMks4FrRdRGakF11y0xyEz2+9xtOOg/t
W66O9wodsEx7s0atNLcRsFxA+CErHOQKA6acn25+sS219o4dmlhBwyYMmU4N6IVXNX7D8fS1qG6r
wCjEki0y12SRHBB+TFMNT8b1GTRtjXqWsqx5NKmOWChrlfEuWT0ozcgWppMzyJVhjK5cBqmtT3wY
JiiPQXDwqsY1PMuRvAAQYaVClqvDmZ8wGGLjY4bMy40kaPTtsu2zvNU+IXiurwk+aknWFL/KkTlr
pt+Hm8nEtk8qhuNhMLeZ2w6S+Omz11RPUAigeG60/P9BNtyYqcOFATm2naeRZudoJ6UtPhLqNqD8
l77zuK7LZICI7Y9B839TuX72aenuvvynxMhowDqBc+oW9TxwFAJFrwzti6xQKC9Z3krLw9RFCf2A
qANE3XMxrwZojEFQrs4rccZJRNXaN6M/cvSPf5HZQFlZOcyWxBOvdkjeNdUnhKu6nHy/mHbQhGqV
Cr5rIWeQrVgFunDZNbQu1fyCAno1+vFmSgBayQ/x8zysIpxiGAzzjQS3zX8wRBFLzjEfrYmk+73G
Cl9vxoXINlv66DkQdGg2E0UwGlzHvvyy1DxVaRpIYSsyVH3p+BldGKO0m47xkPCLEAhbvxoODjo1
1L7y8OfW1bEMfdvz0jldUCO5aBFZMqahCXuqzytrers1yLkEIoFfyWmMHOBl3lei7aSYStR78hmI
2eqi9kYoMW1+XEfYmzNKCZd1XLF7w6MkSwt2pdUGtIs43jtFGT24zsqDGFWwnf/fsdnTyJDnx9q9
BS9ZnWhfFpHrm5IxlE6kWo+xfTacLJPSA1+RI7S4/xCNb+mwKy+d23SMJwdFEyKMAman4AlbiavR
Ru1/U+ASMzjbmTHB6y9pQvfBoWRBc++xDe1fhNa6btAlpTfVRP/ZApDNjAZ653otz17vE9vCgHtY
Gbw3MtzzX38BTZHCvTBcS5M2EQi/zI25WAqLOmV351U0MUp/XJxzGbqYeyRgNtDIoGycLAEfyuXh
HcBfHhGjddnU5XXHF8zLo71BNhKIxj4AeHle1zdePU+Khw6mXdxwoCCp4KRzKyFAf+Yy+zmiGYNn
K0ckm8xVY30MGrgCg4o1cKVQ2pv9YEtuMqPfpq0GWt8oRwZQiAy2FuLOtLreVVcH/f8Rys7l/WaD
k//zJV6nIM0gJyqZxT8vDyo0UHAWRhguZzACizFNukumBGVL4O4819TstEZTmvkC4q2t8U3ce6Nr
7HDDhS+TcUPhrkdZV2q/WG26XuYKBKt0H6ezE5g24exVkX2xxZRQV2p/4JhaQlmFywSWCF1DA7rL
Q77ZbOw6Z2hmtXpyto+vNdGdto2msCivQJS6k5HNuouxOGABvz6pMeZbBF9UzIGdpv8tqKmfrX/Z
VRw6GZnIbJpjqMIuGqalkCFnFk0CDQAsF3IfLk3gFnZfHibXP9IJrOKzdx7QOUojbVUpvy7R2XEG
4vwMuQj4XAUIzGrxU66BIULgS0E94k96C8EYn4BF921s4iSdXRanyohOwHnpEljzOkK09A7mxwzO
ucZqrOWVgn0hZJr69PFOkEbUZXdwOIeI8A7mlBQKO2B6DkRc95AfM7rkU31btsd5KfcZ3exK9Qo/
JIqTacLzhq7HaF46MQqq84LSCyC5boTpFWwTXoHSv3GkP6n587/N3MRJtuMpdly0z7hwKtrCwbZu
L14wvft36ItRWBKEoqq34BmWXd2NlFq366qiOFWFmd7D+iqXI8LzotuHYs5TQ6TdE19NpaitmmS8
f/PlndQzpXJRz2vGacunqS0JO5L1LU8lxXvhaLjJ8Zq/9nrAxyeCXRCVG/QP2WlTD5iW2gRfP3ac
C+X+6lKvwzaYGvRjFUvruMju6zuHLhSokljDdVJNHxEMujY2rwkxOC5hcgwebNxX1r99WJggQdFn
pBzA/+O8tbT0/zNgbs4hJeRlXNR1dGJLkzKi6OmkpTT1qUJVtFYXpc21D45NUusoz7bKgp6vEkAc
wc5xvK/m7oUjkrQoE0htpBSvIUmgGmQ8xohAIR4VQOk4uCXnwhcwB71kMYRJJ+DvS23EKBPMT6va
hbxpXlULVQQ/KK33LDAnnQ+NmRQNw0SDxhCU17XjzUpyebr8KHoboUATFXctIBJd+hs3nkEJs8zJ
NcIQGCebEBJBKTwhfiRnxhZUWOAUHfGDSVpt4Plm5I4Ar/3Zjsei30T8+khn6Uswoi5JByhp/7SB
17vPp6Xsz81s6H5JHmly2ZxJuDDG0N0PLJooVDqGu0U12aUuIghjl8oXkOFLa8+Z0OrWJtm7cMP3
Ec9vVFZPJafCxWdfNYQY5Zzmv24x1KM55FEF9rrjnB20imnZYEj2pQISQ76jgG6SvQM2GqJv6qqa
pR98R1wBAi3RcdgNRRKVksKug2COtTr3uHaZYm6no2yeB8TT8u6fV6QY7owlg/zmnUW8YkjU6QnW
0CPpSYnCQkxgqWj9hGJmnPAiwGFbqhYCpljyR66rOvn5i/UL3Rgtz9Ctku/gayL2DBVTXYHa9B9L
/XuGZboGthIUvBdfuH2NCWh0nBw6LAzW521jQm7a2q+5Y6thYoY0AU0i5mGUGBbQ07OqdNwHMLSH
ZNmG6k3RyeE0KTrlsRXu0LNO3l187g45BtwfqKaR/S4oXBTd06gU0419oYaP5BwIeD3bowMsgiRC
5/Mvh+BXIvkhvyRlyyW1knu41uGoXoiLSK1Vt9g/sxoJ8TgRv0ihlOZSQWKMCcTKrR5ivO6Tg2pr
f18evwb/1g9Y3MzyLReqnrv9V6EdVpOoP88mSKUEm/ZMTaCnXNDMtuV1D9oPpGTvU8RC1tWsBp4X
Zvbg2w90vdDEYesSvMQNVZBz11Z0m3l9gkpI+Kk41PWzb+zYimBMwVrk2meG2JPbLtkKO00tc2fI
uIUoRFME/cbLRDLMTLoQf8h0sG5l9W80Kzq87/um8OYdGkpbT+XEDZmi/62RGvmPAf9Oq10TDlLU
KtMZu81L4Nk5Fkw0ieZZn/TAxigOl9bixiDSrKqZO61FuoIzpsKIE7aoyJKjbmuvHuq1ctWHIzJU
OWTsnbKLduBwZ3AXk2xLWGOscwiEFoIOj4OCBUtetID7nDELFPG0XFQhRlq6ShUUfWn6nssOkku5
ccNhVqN1QpE1dHjHDg1niY/x8pS9M+UoP023TSeev8ZPhgI2Mzng2PtFzsXfEWCrHnN+sXdUQIAv
bzlT1uvua6PpXjj/+4g4qZUhmcZqWDUhZ1bOTGMQ7rBSnKJEDNBE/zB2Gb58I9ms+mXoVFo/2uA5
zkkPpq7ju7tdNV9VuzUNhm0xBdCcK7iI98lOeoaQb9jm482Fjndm8sq17jIOfaTRxRCdGOeVjtQO
vuDQPD+qPrWgut+7LTUVQytehp2j40YaVflKtyXHnzbkPspTHNLODHXF5FbIntQvTStbmDuvbC0G
nMOONCWIyWo0VG5PpnloMZKvhfc7ElQ8sgsmNwT/0FKHzNet9qiUILyyHhQpBf+qPyPoLOPhk5XD
crqstOgsaMwxayblExCSFAsZr5jsdtFnqlI0o6oILPExtAV17Djz3axQEZQ9/BI6X7P96WCWmxdJ
vdNy0i+LIELhrXuhIAP/G9gEYy1+Pfk5W8T7gyQhEm8NUhv25pIBsyRcElORtoGN5npWUvyYYrld
dgzDBIfnA4QKhaDmI0zW3Q+jfQS7PCmuKJ6uvRoP08FR7U5EhvNvULe7TsFgIOwyDjeFu3SVTFFS
IxfXGEnFef15MCWbuC4zEyyT7G3iyvyXIaVog7qRnfdI/4sTwbSix7YQfxeMUoPH4Z53xKD2Jajq
rcGZ4aj4bWrpckKL6l38a1FJLMXMctaf4iGPZBRwYTfARUOrh/3rACwy3t3bhFBCNzJzFIgedniw
XMryWNwqOtBTvWpPGXLwRWdVpweZbf0yYQwzsUPtmHTzgtbipdHadc2T7fSz/8ixD5g4qfy4PBoZ
+7riwc6rZ+xkdat3iN9N1tWwd0N9BefQF/l0Hi0lZa1lqRSdJ9AFO2JlMvmeddPnisCZRjWqDs+x
aPmaESZcWoNQGJMRE5bIAxtnS14zWmTw/PqrYDUq1EebzYQ7xHkQT0GLKIfozyHB2pQ/9TM99YID
dlkqYkyZJqiaveXxKt90U4cWlYe8jagIbj87hzOkocYO3KWRWODuOKompQo4GWJGDx8fm4PDOEm8
WrZXUdypFkxn6spnT87F6LxNYbw3yFPg7+4LbLG1SChaCvxVrGDqrEa1r9mMvQr92bq8WFTLe3ig
q7+NRCUheL2JNaJ+sB6NGt1cG56kA7MtRHffbegOGuEZzFOFT3zUvTvTXqZub/O2UgiFGb+xfF1s
R7IPunCu00oJPNskPHgiuNt7P1cC/VWP86nNARRis8ZFaS+/BielPfd5qt+x0SVTs4prGuwqWEkP
rwMggReVNXMNU4VcSAEixthsSWRurm9Q4wkzdTvlOMZqem72Ayr3E4fXoP5U549lPmtgF3e0Gdb8
FrLeGbjrZCyJIOat0lU2Av30a26Whj3312i7YSluYLEhiOvXIpS2E6qZc8RrZ4zZX3TY6NNUbUG1
1K4B92H/XpA+o0YC4WZ3Ts1RkLJg/YCmChvcg/NKOQ7FxOveOqwDBojM3fhMVR5x4nlXLL1VIm0x
FyBepoz3qIiXEWCmw1oYSYCrpL7uerDjXMOg2teBsnuSyGWFcaUNT9hC5ZNtTyAj41e7nZhJgL7R
3B1d8hTCf7FS9avXiwaMXxzkyMjV51Ar0G898jW4ozSRgvudm9fXIfeLfOIRmzMHjk1t3zKlz3gS
9fuWYG/ELQgOV84JxeKZEuWqO5GV4Llc2tF6y3MnJIHmlgmgIIlfq+T4MmtYDpMSXzRhtEOJSgR4
c1YtV8K5/dYGdUpgpmdfF2/QV5aV/fXmPkBF1CsYcQuYDg4H51MOKHPn4eWFxoskVKnc1XLbc131
fTuDQPBIxqnkLYidQNju6k3NuXrH2IobpcavMYLGFTeA9ekAdqtxGE6dVfd1IuKSPAel3mDB7Yny
HIInZh+xQWHHoMOeSnnfHav9U2Xbv0PVteVqf2TARfRSMT66XJpjTnzT/BKA2m7P5eyRPoYYtj14
FHQsLRiaPhgJMIZQMJmAHWvo5KTnzSLpf7naKb/GuqYVMmDsxSY/pXSkpL9vujErTpzDng197+tP
4puDpr3RaBkHEtz3LFtoq7x4WkRYf6uIH2BcSPCptLJc7XGteQ0Ogyhi8ZLNUNDjqc7uUi+l+g4G
olbHxlsNH9OxfaYMMbMzzs8nNt1yIihG3Sm+ATYAOaDwyaLCR2MZXbnU2XDNskxRaoybbN6JoI0H
UxttOcuiy0s5lKB+RNNEJphXOJOm7DwB9CNGxsxucADtAgl8tAW1q7WYmwdYsJvVCFMEoR+LmGwr
BhT8CIAOyQV0EBrZlOD6WQRuExmPWChI8TtPwcYQOm9rfgvf2Qp+VU/jZFeZYqGzyQflLiqq1paO
jQWIvW0BDvRXNxfStNl7Wg3QwvBV12/iuarLqiUe2D+vHtG2EODHmYgMKZFJw5XTJ3jzNtU+iWB/
rOS5a/qA6GH6+KBAdtytZoIq3/ro9lg6o3m0NVOAlgjIR0gCJSMvwiyMiUV+nh+5zweucXbNscar
zjdAef/j9fmr9wiKia9HF0Mw305MEE1n7ua++tl21cWqYJ2ONs7cd1iz3Xi8rO4OG9jHsXoAe+lL
//b59nuAHITsXLjFB/6WoJf6MMB+elmlkkeZ2coRHwFw2vnIETH66HElLTxCaKWdHqOjjj629QPx
ZOk5eK1D29s/VWMXncw5b6fp1UGJALBGGC36c3DV/yHosSEnNfH+HBrEQbvEngbX0gplrjc9SnMi
h7X2uhBSMuwVR0Evbe8Do9prozhqmvWIWS5mqUdaDa+bbiD5VEerIzaZZqdENpxDohXoPA/wVHbO
jwKRvE15woJS2BhpucjdmdGfhBL4cHTiJACxpkUDNTN9fsehO5gju9eW+vE+0chi8L2UMSPoyQGW
1RZh1OKOBjJ5p+0zdJjkH7zfhUWD8FcfgRHui3oELYwHpyckdeQSqyyMxwQTSXoqiF6DYosgbRDM
aQO2kucclChvaYgM2iC/PN5Bz34Gs9/ZNWa4Afj6/RemW9bj6lHUNyadLOAr5ae2387G4R2dgP0H
Dpr05tcx9hk9Ov4wdzBXanp5WD3HoY9oq77qS4USucTJPdogAaTjjQCI1EF27ngf4D6QPFR7uhcw
4AINxQn2jVH3XxjLpuuvk3xSoLRJ2xWMp052h2rWM6B6lrROz4DUs5v2mrA0ZcFGe1VZjDkY7aZw
Clw9bArp3GaX+0VB3FrmIjiwEoCtVD/cytuzTqDcy5BD9pzn5wCkAIdkvCmU3heue0bsNa+BqdiV
rnK04SN4yrLZrjj6iHEH6Q3mJQb6cJw7FUYTa6td0CDtjeHB9d++Q4Czih24zDdgHSuTTVEu5sxU
hKKQRj6qiWFzaAK298LhUTbzG0vjCyGpEq0JiPKc/zuvGPC5Rfx3vDHEd46UYO63qvkyN+habVze
G7gG4KdnX3elwAITPVYFZQHC1XZ49QVDESmoHPsdt0feDCmkS24PJrqY8h7Be8VzihFVOk2ZiI6t
19/q0wAQOXH61FDV7+yDwMDyTIFm2WThTpR1GK3ceJ0rfpsJp8213aeb7qVP7sICyZGy7lZQsZHR
myitZuPi+zTGteu9bDobFTyYXqpqyS4Z7JIKKLKbFhbhdLDD4xt827gvErunjUeLb98Q3Xx5FvxV
Xi43uMYjjSADpGKz4kGw7EkgCAK8kOr4u3NlXkHHZ2cqzgfUJd0FixliLX+bpyoQBNzLCR3kZiYi
2POhRKr5NKmH+PBdswo9V1gG5EhqBA/X92zeJST+bpIxGGwnjbTvmo0PY5Uc9HLN3gDywlaLhuJI
P/pllfKQ4/vfogyxkN0WIKez9Tj3bApA9IezpalMgqE6KmhZUpsQ964eSDLhVTNJu9KXkG3wXmwY
HT48HE6hQ45gmsYxS1EMzX2ucVcYfrWCpLrRqIcNDpg9gHT3C/6TX5DJQ04bKudKASlz2YdL407B
U50KQq8fYZRpnBgB4sHdbvEzuxZK6DXPUZ+CXOUd7AzN/DLxYV3IcNhSnDrhVV6cysst/X4zSJ3S
sCMkbztJx3x97C5V057hrW4IKxHZkGUOM3fhMi/UDGY87NYmvSeXpaRwHECWurqzCoZqZNNFd70D
OvsRH3sGqxctVbUF/6qSm5rQOqkwNlXCWfLEzy665Iad1t6hMvFrwGaOr7SyjmbSlAWejbXNDlXh
8VAt4bp5FA6JF/3QRXV1uxPYMeWvEYzCoaJJieGIj0Spw9vdnQzv7STrn1HIKJAfFQyJegtwNIRM
wwP4tCo1bJsmmgqI5KSW5h9VsvO35/9Hv5sHVHcYKCBVeW4y+ORHUx7G6Pf8vhw7NE0Pr5cazZl2
iM/6Du4dHpECY9z7rrrG+oLj+c9uijd8TzVgUz6lNtjXIdVROCYElFmF+s38sC/nGFyZcrCpsMug
pn2sj1gs9ZHWLC2H7Rsbx7saZw/e8k0vI7YnFf4iBuAR4kymX5OjVSFMIs1eeqdXDptu5TPSfxYS
sWJ+lugC416hZx6uhhG1W9clJV1DSZq7MMmYQ4eWuS6zH2OWuRl9y/WLsq3nbUtjUrUgoZnLmHCj
0XoE7VBI/xKnxG6mvqcgA2+yTDOdXKJDzP/BeJhnN118bkeUTQa49i9il9+t30iz9+tDMXD1y4Iz
hNFvP0U6A1lXPhsugM2mRiHA4fRa8RlwbZkrnSe8V7eqXtUUS/EFcxE9PJHfXEatKIzJdqXMz8IG
oxhYaTMTICKMRux3DV9wkQ9n1H6geukAmsxGnC3/uZzjRGuLnOLboVDGALIY6FiJ/o5M5zoWiDFz
fLQVPVjtT6s3Xe1HqWJszFQgGw7euaY8tRWizYuVBB8nUcNWSfN0etLrOAHgJm1gCYWqZXd2nD5D
tHn4JfQHMFnJji4JxwjK85/e6b7/z/OnafQCcmbpX0tAXQ0+m3uB60HAFXIs5meXYQt8Hu/+d5fk
IoAYmaT5OLLdDmQ6z5uU2KBLEkhGfHrfxfTFrMGajpGXkvKh1YCv2Q4uh6X4yIb+IGB6qV8bmC+E
CJ0+DUpRJau+yrgNnPWyFE1RNRNL0eaCvJX5FkXLn/rHiJXqWaAsswE2Hi4VNtBA2IgwnSQEJuzk
uNpvY8HWnELADWXWivFNIszxBcAX8WuLD+/ORrQ8VQssuKiWBqZoLCaoS1hkVHyU1qDdv+icM+ii
YzlWGuXnJTTD8Evbrmr8kiPIFASm5QOaAV/eDja4vf6i45TveL1SEzGGbzs4iihwseWTpPLMKTGg
9utM7eaDmPBdAaVTCk9Tv2p5+Fk7fled8c1W7JhDay5DyU1lnY6TRSAkWWrnldvOmm3tdJYLc75u
nPDWZ65XlQlB7w/5fqhhLibRv+hU72pJ0SJH8AKTP6UUI7wcoiBeWojNIfRfDO6AmZif/qr+e3Iu
wAAFj2UQvMNDgxz1sSw11LSD1X2Lvvn+auWvUWrm7PtRoiKTpdq9AAHz2G4HyEu55URr8pxmKACs
1qMpnX3Kqs7P5SOoJY2aeiW6tv8EIcOF8aCeOt20miv/8/OGiBjf8+jLvV2+icUUiCecMiQ+8e2G
Hey6o3nF/+26LSuRwpkIZbU9tUXOAx5XI+WDEu4EQk8jBGcxDGm6Bw43jEMZbC3qsQ5ysVrLrqtk
6/pK+M8Op5pBx8BkqUG7ZDxAOhqbRBcv6VIIQyVNuvDWYEH8l1ZMWdZZRe2yyAa0Yq2GAlAbb4PP
CaLkdNT+XGK1BeF2Ru1BRLNArx+Q0eJr4CNCd+SAWfFXidSt3W9gdcNObjqgDmSDwUM5jSdjP8kV
v6oG9N3dMBbz17ojSEPkqDy4vT/svMMZMHOuP9V5DICiZFFLPNuIdxQL/8intd7Rx4evHN7uW+5r
hNchwgVQ+/U4bi15V11pL3To2R0TlJFIZ907RNrJp8hK4IiinpBx49EN79Ox8W4Xfvxj9z4E+NNT
ZsvP6l93rBBKnLt3DI537wSU2arW3isGmEweIkwhCgmEdMa/SaFO2/AB3f/tVovHgr1X6RVtmz+W
XXcRtYX1WISggzL9XU8K0VHZrLbGkFH26mfiFja4mM1aXLd3MgrNdoX8RIbnQPhXb0On+sDQgLov
s4bG9dj9CNffhobTS6dZJmUAita0eudIyzln88MOzXVqtC52Vy3a4XFJWIxDtD7Lj5QmOrxeMdFH
4DLCNtqw/k56DZJ8gm0vsXTT0TIUyPKMgPJdGR4GSbtdFPCFYTo4CGEiGA8Q+KH/tzX0wCe9lX9Y
YknmBSpz8+t3fROhN5lsg5YGdKafq8o083UHvyUhaK6XafkgVRCMIqUh2JZnks/4kzCROJWZAcPv
UdrO4TQNFOIahphNz02gqzTKVXSQR1hse5tUXs6AeR0SGO6bGoJP9wE4a6oSns+Qj4tFKazBNbk4
/cqO+/YIjABJTL0+7JD5WPta++rGCurjP+yE5DcV+4PtZJ2Z2+YKjViNLLWjmvRk7ayRqPLBJOvx
TJrAFTPw+W587BrkCNOJ43qHRzH7bR76LE10+pbRQFGbRi2Nv2Wtf492erf/ULepkV6PuBwNYg2V
FzLyOXxV2puEB461wuJUNtyPouS4gKNrTMmRsK1X3CxcicHFhXk0uvwkX0fjC6T9PQo+7qcChRsb
Q5EAQeGa2LFlqd1SS49DaV28TiIn8wiJ103dN5YHCTU3SVzFuiQPBz8gV8DOtoiS5Jp3k1+NEvG5
hXxrge5aKt0RgUvwhG67TKSk7O7VzHZb6SgF4cXFlEZBglfO/lG66tAhcDZ8kWw+hd+Y6AK8WHCb
o5c0VW2rvPObY1kMO+0RIhxUlVZ1WkF0+XilxIfPpNfx3CTT/kmq5cjgDtJTO5nQ5wMX6Emt4VXR
i7CkVUr+ATng/60PPb0KqSHVQjQ8P4fQzZEdYIRDbNf8EJ5w2r+goDrNmfCq/hM0WmSFcBWtHFje
9Jg0fTd9aJrlYHOWmFb6vLYDcpW/4StBozDjyOEnMYvO3HVai1y/UFJMmvIAX5k2BfX6yGNUhq5z
qb1mrMqLwwqzPYYJx2x/oQvO0RpujXMjLVAIQbfRS/VkeX+6kKS942QFonfFKxZLc149/nvBpab8
OOcaNt3/hBpd+Emqisjb4D7zup39Vp+axKiThcxKB3DfBunROyAPTBf/U3IeoMmbM4v3IPFYCwjm
PHw0Pt4AhiZwCljmzkeydKPyNhUbHdCTl/iBDA7LDmNgrzmULbJ+OTfUcj+Aa+zBLoVAhXg5Lz5i
OaZXSBVrSmcR1lhcO3d7J8yuFd9jZ8AlqvlpwXqv0L5Vw0GuMcgg0L8WXhT+q/uACUPurn18lvI9
r+XLsdk61vkyAZulPS8t3u8Z1dILMkJrscOr+S5p2f4Op0JikFkEm6BWQBF0dRNP95nckYG3rd8M
R5O8QBF2juhgmCz12cE1QG64JAkx8HPmcRT8JzGtucMDk3oBQweiMlvSv0LGOprpLoqbiqrRicyY
N75DSB+Wa7DgmXqnwz4egjOAkuEOoGcgJscGjqaqlHtrc8PzW1QQEhvwR6oPKpMyWcSI6YwIB17Z
pgsaRwT38hTy4EDKkHgTEPd7QgBpX037xOzA7VWnl1JIie4EZ+keNj/HkVD5XX0C1v3+Byld3VCT
e5eG993DFtXLwAOxHvBVJBd0o536fSLdKn/VuDeL4O0lr/7GycSl4d41zyateJ9ze8pdfq3nT1la
oJZyN+8+Ljr6MneZl+KDCI+dfGe8zO5WiHbyeQWwvt9PSEQFq7V3kEXbVrcDm37FmG0IfSrgB42+
dzvMJSddMnNGivJlh1v9kOdcPnuk2ol18P6WcgCFamfweO4NzNx1DCHe5owxXduiO9uMbede5SEf
BBQx2XTslueXPpM+VG6ZrQUCwG+OlafluKWxetAhnpZeHv72pnUM+F7BYd5B13oWRsPyP16U9TTY
ILvY8P/PZsGFcGjnIrmao0ZALWu05ZNGXCsQ361KxtZoHarXh1/f+2A6ReFxxLEn8fsQEp7vh2p1
A0qOT6gcZ4TrrqsW+ocIXDxLDta36LioaW6oYow4pcHmOkFMpK6Kvhv32bV+gy402JsF9bWQ5kd9
GXd9PrK3VG3EZtxTy47p/wsM2kDu9QnQuXrSk5OMyZhhtTw5fl6477aGXWm4ZjYs8uu8rh5OkI7n
GmGOP3LMSoHfQ3Lyxrw2LWo4jq04wN5JPjh/aJhvBDnd3470zrg7ulM5Xx/QM7gxAcoxqEwhCN3e
jFVymuHgYgiZx6rBmn3cCllGRifCCIAboqxDofMRMwVvr0in+jhpNYNMKzqwIYlNHcRUZN74Dx/d
LPz5ownwWZFr53jlvOkSSUVpUM0RormUDadPcSvXMhH+h4Z3Q2aV9SAubLrdwZmN1OOkHQDdKDTu
qq2+If23LZG6zCBeMnaLR/ccm8qIM3uI8gPs6rbfYtE44ImFpDcosfPUVQHps96Ia61HlRhQ6r1n
jYOtYy73O0Dlyu/s/uxhqnytYcIkS4OGDpDzhBFWq1p/uIqMvIbCrdlc5UYaPtQJ77b0rP8OTFZC
T7Lw7gtZ/bw0LJY6iDgHIWLSJUwDaexCtIzd171GftuRQ3adx2tmT3IERFztNo2pNdeaCFSyX+TT
cpjztt678JsMUO0ip03RXeOREU76w0JPtJEhXnrU+/wBXu6wq76ax3J1pKjRY3ovZMRr07QSYjw5
WpG9QqbtrohQ/DtjoDKVN6nfDN/kJjyNvsRmewMgvx4uy2oqEa/OGIAoAqBPxWf4+lYLKM5tqqMr
hiLnabGqMN6oa4uD67zxEcGbbcr3uiRrqEbPplE33lA1BCopulK2NP2xrbv39tyuTB45m0v8g2vz
IoDnjOcPcPP6Rk6U3srl5p+2FqXQ0nAiC95/3Jq8EPW3O1hLPPnQRUdnnl0RuXjN4JCYPssobd16
L2CmaCkRD+ijRKyWDTWTp1V60RLngVrElnlHL98aTaZerY6sg/It9QO7dM5BvKJIx57FggDQox0i
9YaQcWIttlrnzCuX5eCqZEhNQGFujzzXiIsY+8tCPyNxCkc3bzEtoh7YK1GGC9lQAziffIV1e/7r
yvBJZj4uaW/I1iXOt7iLmfRCEEhj3f+elXuhyXL8b8rp3YbQyX1YhPaQ2qRNyvYfMmWDy/vCjcQD
cFA6m6TAbuS5Mfb7E/fMIm4h+M2prVrFh9F2VCx8k8jP17QGVNFRlDiSdV2Ufi8fZWUUeU+XGR32
jfVb7hA124mxmCzPgrpZsQ4buR4drYuGHlNVp8fBZIxcoCcHU0C48rhFgalQlMq8tB5LBoIl1Fbh
5IajVL9umAVJbWlJKtLPzZTZsAlEO1aOsGpapU17axO6efI8K7Ldbx73TpeKZJHs5JS90ajXPZch
cqGw63i4OdpsmSyjrDpjlS9SFJa1g9T0e/5597JQGoG9+7NvU4QsXT7NqxfJwau2VTxR+NkNzDj4
NfFWqZss1IrfaYxaHMkMzR0P3Fw50jedzvTLFH7VWgYZQfb5jQIXPiHh9lgPIPnGBuKj0M8a2wKT
b2rTYnXpx71vp9ukLbpXxrkw9f0kCeS0GsGzbivz+qsAXrf9WJRvq/mBuLG35yDaqmzPTQJT1Yf6
O8L/wcYO8A70/8TGmpXBJ/3MRUmX37reYLwjrwM3+vuL7O801zwOMvPV8uw1HsxvbT25KJp1LeLP
uNNynws9wiKFtBT/ewVY6qFF2u+c+UdE314H6r04qqUjWpBdx6tG1H8iZkwmDU85OoaNePjI82sG
Px8MMKGI1ox275mV8J+3pPv07YmKSyCVXSjU8bmUcwJ2N4FA8kwW2kta3lu1RJWduU1mLf3lLW5h
myWBbI6tKURVo53L/WT8zcymHuNCTNqALKqQN9Fksr/cBGKIFNGprDHWWBfqeabOuf4oVXfETBxv
Pts1ZqjPSmEgdlO9cNr4zc4vugoq1VHtM+q4pNgKo2R7DKHsMgLf4Tv05geWAL+kN2F2oGDbqGoZ
E4oWDmCtnTDEQWwKUHf2TKYT//YHGSmvWk/6IYhdJ8Bel8zfQSo0skd3D5L0ZZXm7IMECtXVgU6i
i9G5zRrtu8wKioYzXbXFqpZc+h7VxdOPjN4xx6GnNyqN/CAZD9JJG9wfFnTtN1OdRjZTSEzrtZ8+
xHGeD9pBjANlD0jyRlzEyFmXJZe99v3NVYzNmBhCh48vpyyDrQId0rEUaimX4x67aakVLruPrO1E
+96dxaBCmAtJM/y7Y++b3vFfbqcov4MeAZpD6WzRE7mP4xVrLvVMBwzeCcCtay3sEmP9MRNG2Oqo
f+c4BfwXD8H4uCeEKDYd5HChHlNIMALEqiQakzJd0jy8m3/8BT/ntpj69aJ0uf7eGe9mgQKmMKi/
BGvYj0tPqHuMQO0yEiyLi4UQlWTK2dZ8pfF8YrLLA8/cUMR2rFCfEVp6pHEGu7Qft2Pg0T7S7+B9
261KqJiUg1eweAkG81Tmb8UdF6LVnRpkWzU1iR4iHfSmbBAiiWbba/LN4rEMxkI+pZmXwLQ8j+an
9EoQclmcoCCLJaHcrL14og3R1rJCAXq48jC7wU3dh177H067Vz840c62KHqWw43ThT0UmFuNoYZM
WIho19L1ztVibxWUElq8Iu9FDbEiX6Qd9dz4TPyfF/RmUAicqsZlwZ7E7H0nHTfDXRYiSSLEjcMS
P3gt067OWEXthxppjmURR2DxcV/vpBe27QWq6SeHkLeGPrz9b/y6wKiU9ETBXEVCYk81rEBp+SH9
/95voKYV9IyuD6w2We3Su0diH8FepfT6JyMPU3M0pMeBB7hgaFUbXnUOP45Iie6Aqix2Vk7ATTDz
ihvnRwoVqyf2UaqmFO5ezAd3yecGTNtTlA9Lg+eRAFxY5UeM8LJwTm6+OaLhXb15iowK83Y/NmBS
Jrg2eHTDgN+Lc6CGbl+gB2j2WbCrwqvNtKnPRlWO14d96+fEJTqPtsC9cWOP+ZLBzQ6etIdK3qCS
uS3hDflnw/OHEKaGT6AEHkhqh2bEcquPxbCEESXDoeJFcxcF+nHOtnwTp3cScY/AKoZDaDXRPH1I
+3AkOF2bLt+zrPIauFUxt4wBOZlDbjw/Et08fngBhyJW3dlC2yiVZxY7ohf6T7KHDZ1r55GdiUZZ
05+kfhDN9e8ObJ9+IUHL7BzvXOw+4TFG5vej800OY9v7tK6CnkIzAZVYZNHyZLO9tUmAhtbY/mwS
tYhqodH7zHpFDH3r407nnsraRfWBQHB475frBbn3G5FYW9ndP4rsuzOA3ImrnXt1CwDChQj192Tq
/PftK+B+bEMaiVIz0btYAxhGnfCfH/ax+imJaIjsM1sWPwlMFoMloNQhlJqycwzUOMY0WHDsutQG
2t6v/ExAq/+uE8jJBI74XRCg9QhAl37SL3IZl0qaGRXiMAzxgc3rBzWn0qwTcHuTRv87jZEG+o7H
abvYSXKteatzSdmW6lnTDE89yWt1nwlWhrT8jGP/WQwgFVE1rVPAMUz8o1fKwOtKoTCgMjNaZDxB
BjoVnGV5HMGcWRyI6mcuCv3fQWOj09F1kJpuQvSST/rWrIT9QKmZFpK5IvKAXNmQlJJtBaCLNsLn
zysmGYUJTLijszENVKe1qqkOhr5zCZeEz1qSgb9O8MUcdl+d+Gp+gpNIR+BOkpTdhRkEQF/jSXa3
0t9iz3Wqebu//SRaGoEep5qyuUcLYd2gunOQ3jVrOOmOj1RAj0zhMPshCHTBPvbMV3et+VRJPe/O
ZCfqVdCiVqF+Wwpwl+DHmWueXYBr6FinfAx4ejIdxo+tyg9OZN8hsBVyLNujcU6HMKWI9mfWfdHH
EF+Xh+G6TW+RtbfMILmrUCalqopUHDpaUQTtsmj8asNuZ4SvJBsGt7tpU8e188ID8CuWqgByZrQd
5jVEOZdu7v/oCVXzne/XCofW+bNofz9ChqH9DMxhDVhjjxn06WsgLm4CKapWHb7IoaaipZndK2uM
J94I1FrfQCKtDkrn87fJPihZnAMs2rmc7DmWMMgQHhWgCiQbf+W7b4gv3oZsU5ZzLC/ZF87nmWVO
SCMhrXIbPlRsdDrOjbmMXeMH7OIJuVfmJT6KjzsAtxEjyQbwt49apHoc8rDMzbh21kQhE2JRFjQS
D5selP2rhDv8h81q+Wj9MTP6fzhPGmuhx0sNm1nttVR2YVpalbQe/ySStV/bos+ZGRuBp/sX0pdb
SntJQfk4yHNXw0ffbUN/fScZJTbblfzhXuMTAdMfJqrMZQF4qx7x4JU0MSYIINnG5G9lmpJO0Gri
JbBVyiccitcHvQIvUPeyVZzdV3RlEvpVyKCRjCXymNdqoCDEsROtvKUOedsvGjxygMEQJrvvlIrN
S+ZZ/P8cspYVxEAnqV6CB3Mc+IA0W2pwzurM08vhlVNZ5l9M9LFSwhk3H9C551QmdzSQWUFSTcs2
rgJmt60MWj1pZARgJ5Skdb8FkOr6JfG+q7GhckBEMcsRoUDrB+843zuBGyukY/n+SpIeeJcgrWeZ
mTF0FIOqJfsGhDbyuUQNBJm4J5SO38CqIla0ke52JVuOMn9APtyJpO1HrcQsba6MifReUUIgjEZo
NKTbQM+Itg3VHH9AHRSReTYnrm4oTI7j79J9tJVIkoYLVvIThdsB3ITarVvY5K9ur/qI/+WfF5yQ
9esGnVQkeeSj5vR8e2lnb08/FdR1DJvypvbSxxcnv6V/Z2zipXLJif+JCVFZS6Ve8EWP/KjbRNLB
U6xBPI2z/T9EjQcbMFdxRevuIKZxNFyOwT2CP0t0nZeaTqufnAfKlFuVBcbMVUXd9sH0bO96wMPv
kPSN+FDH4+lvxeRLwGwbl1jwzbJvJG0YLdcVEprJMiT8s8VHZs/oRldhJaGpdKKE32hRxmu9/rwe
h/4Jqzp4evlwMOyzjUUH1mRyGhefEz1XjkERa79L7ppXoUy6vLcsasctSSfVZ9pBGCs4EytWnXsn
kZOKnl88NkxRLjK9/fJQWubfdWL/uOymxiXilNDGOkHGEtt5zhu008LhatCzosGBbM6nJOrfEF/l
pX6OX3ms7BS8FjgfcTpiVG+4ED4u+UKWKzs0XDfCMSBdAGQcmysUcZc1c+cFlK3zY7tnHPvzwyML
1dIJ5CxQJ3AsuB5WqjrzbSmbRtIVMCAgrbnFRw4mUaNEmrmrvxYO1gnsOu1gf9APO7mWb6r3VGvN
RGPaI+svIrQwlKTsxht04vt9hNh5gIArEsCipw9wed05i2pQSlNYwwqhBI2mMUpRj5AIt4UyrlrB
9QWbs2qaWzJFPjLUHPYWEdKvAQsW+jqTD/pDJMA0fXKgmSp66CJ7fOHViMXo+CgVPZduQhpOC8qL
Fqr/G32i7S0VvBzquNKmXI1icGLOPN+D76C+3NOl851+wxLr+wj5bZhUHQDmjS0WfgPvBi7simv0
iSNrbbYZZ+lodHSEYrS0Bx5osESTwAwafA8VdcWwfuzDa3Asuvwf05x/oMgbKDVjiR3EjHkzHlg5
UO3UpsYFCILuMvfj6iUffGSAnbGVFUAPGwPMeasCqDkaJYYgt8vuXmWSxQStQBtLBgoqm8iTHL1N
StFD7wIv0wQ0w611xcBOo4TON/NAf4i6NAN13SyV0vthMeAH4+DzBr1Wy+zAI7GElEPMJGbLCzEn
N6meCwImPSwStIuZC20ctkDli4YlDrapnbVwpfWU9zeGhNDf4bMttDlyEVd0fO41+h1esmDZgIjd
0vKPD86loXCwQk2ypg9BhDATkP/dukUtgSkxY7VxT621HPDmk1LRIfNxwuFVxPAw7vQ4etHFrHYn
eI5ptcpHiMXZTSRzLEZhrd/ojHxENDxXx7KeqcrV86DIL4cAPeGZOV7LaOk29q0gR7qGTRDHAVo3
EPFFYnBDDnuAH3XteAWw/q2Z0m3bupuYQcLDrfjTK6KcdjdUjK79iNBgV+HFPnkjYb/+Z985wENU
NyqBele7SP8gYJImrLvBTW1cUwAMTUqzLTOuta2NuYFAdsY70ulQ3TVg9g8x1FEs5/7MyzaM9bgX
qEbCrLerjG7XkPu3nHyb7PWbgNn5gJJp1C1DRC4Elq/2sNbdRRpMfomWNtVNBboByqomBcOnIMm2
VTqSBWuhZn9J+bXGfaxp3XFusz11pap8RwzzorsuT9HtEkx8ZZ8skrRwWxL4Yk5i4Wp08iDTHodK
IQ3NuIRgAglOFy2i7Sl0VsxXXvKgNLqRtdbxXrQcsi98D1b3t7uZ2iTxqcWH9LO6pgh7pjfasiWk
oyze0uCglQZgSPU47YlaUFNrRJqAKnHcIM/dG6Z5hCdA79C5/88drln9UpCEYDbwybVcg2JyLbLz
XRpMXKTiz6gH6bzCef9J+LjPjVDPtUfo6gUisdYQMYgw1eMNRtB6riQjplRmw1HRxG+G7gGD1KRf
Lav+CJ6Ui6dPMz5HPb+5YDRCjN9+yTGlPSNdxxSVfIZpm0QUZlrPpESM+3x4CBSfUHGgcJrEnJpR
hRQkTFkvTsqxQjcDgaJkx5I7YyhIzTCZxaKQGW/2/G6XR5n/4iNB5u8EvAWxRaFDGPwfcoeunIFL
i7UyDSvWmx2FiDv56LfAi6h/i+tsboHYPBpktSl2mPjhvUoTNKiddOjzJIB8enyskq6JM5VwK+Hy
oVhkOzZJTTMv2q760cgDFHlRKIyosfytaguUreMXCdKfnaO8+oRDqZ299ejsK70uIwN5iZjvIQ2v
C3y6v+QD7tTOOIw+uRqL+kUrPeV4Bs2mkRxL0LspSaGz1aX3n0VLUM8a9OW159mL+u+muVesnA77
e2KqbA1JYpZ3rgyCRndCHv/7yPv1ew0Sy10GKaLw7RthEWdpfDefsLvCC1TnyQSn0PWT9hxfbQC4
YnJA+UBea4kx8BTugdbRIwK6ohs0XFidjdAuApYdlgAa0/qAAVSy4qFbIdfn1zwHaI6GJ+OSvVnk
IhrPpIhNwAzi3kW1HPU94YZXZIwarUvJuN5Cv4rCJ0Wh6g6+7ueSjbGIn3nP0IzjBiVkAz6PqmKN
qQ5JoUtwsDTgzIkW/HeQ4xaoyM2spDEKshSdVN4M03a9MXDtn4wPtm0mBgb4y6KVT2D5aEoVo86O
1ZM4IFWlza1luQ/tNh0z8rxoHnIMTd2433pGD1WwSikrNkkM5Os1m3tXWoIv5TxEktS+yBaAV0k7
2rlXEGy91wC6z9xWo82ciOr6//M7r4JCwG7CUiEfGjDPuRBzX/PsWdWkGe0r2fSm7/X29+YOlLcj
VY+i3HHcBDUkb/TnndL4mbJP8/7S4s7EgQnShroOY8myzNuaW9iTz7GwYHVe8Pw8dYxVmK7R2kRE
NLB68jMoVis3iWfOyPUBKQ3yVUl8fVo8JbEQk5aRFGKQxhdadypOK/qbXh1zRWNwl0aJTUvAujm9
ZxM9Z3OK4Jvpzphse1Z9ZSYKZuHMtYvEQCLAcO9jx/YK+z+NsS2Rs4rmjzQyMAD4Ix5NnMiXTxix
JYyYvHr1kPcJVek08BB0q1hkQMPVCV6orA0goUiRjeU6q4XXFl87J5OVjL9DE4vHL65PAQ0lULhg
/ZdjfB4tqxQF43sAoBaNOcdjYLH78BENkQrYEQGj5C4h+eAQ2oubpOUYceNEtt8dPyJ4Ul/fN9W3
MVmXFVSn/pZyh/m93Ah0tk1fr6dDQfZZXyI0T4U8tm/qlIUlF7/b8gcMVrIGnDyD0ntxJKTDSjWJ
8zfOL0OuwVbIalWtEIJnPlIfDdlGwOOgwVzeWNxIfTc/48skaPS22ZUGiVdxK9u/VYAzZ74JjGH6
qk7IREWu73SxSeS9KXo+USEtmAzjflFUC7JtWgUEY+Pn/IVCMG/fwZi68NGfE3p8UgWpTONq8Pzl
wsjoI8wZOPo+gppxG0ihASTpy0F57f0aM/kOSNQvA3ZdYEZ7aflgmMoL11WT7wCU3jZ24066T2mm
5MxGNNbqa8XiZKtWhtAbnwx3/naNY+z23w2Y8sKIGWGyTs5q82XTW83CafIFuNR2+suQfDTI1grm
lloMfh0xrQKzHJm11oe2yal8emL4j8oFrTLpzr4zJrJiuw82VmC5f49wnXImjNZq8yKkOqp4pDZK
4hGw/5xKaswp7AqgYf7fwhuZEr0Jg94y5++LRBjoshtXC466QuXL1efzw+hO1qMnZKiNdxPh0NE/
3TgyBH7AAuFP1BqF6WLwLQ9EV2b0BPddk7BH33+LO8eOhI9RM6IkrG2QF6Jr4XGCRH2U4BM3yGsy
faGlF/8WBNBg68lh6TSbmt6YYNcqO5y7gvVG2WfZGTpi4TT4BgLAndA8ZYJMhP9cJTSviDei8mrI
40iDXb5+R2INsOQenkgGR4Wlc79M4oUayKmI4h/oumJrTw+JIoGzxRwdidIgSe+UfVtvvBJeeEvp
Y6YKF2M/Fz26EjdqzxzExBE/jUyWJXUfcbTKcRuadQyu5g+S3FPeh/e0sTMNx+R1Ktw6/SS/kPN6
gONQixaqEcxRx9t0KtZLjoPJMx9lntExsSb09LbLjQaTfWwdbWuweaLTO/Egq+b+ngaQl8Uz2cro
W0DXsjojletqADTLBK5ub1tPK5jREdcERRxs3K/4p1EbCO/dlxVHxrgr5TlvUtycIxjHc5bUOTkJ
UoW3h40DWQ6JbGcrxc12SxqMxTlgYCj8GdrslgSk8FDjuYHNnFoLpO5GTIlJDyf8yA1DaiPowfg7
RGiyHPh31+c+XFH9nNinAnyqvR3KjJ4iRTY+A7VHWsuK7AhNu7rUoaKA/+sl/g5fC6UcyHz5cZg0
LxkhOlcfFbpRK172He98utAxBYt8oy/DOtik7MSG61LPsL93xcKr1GTz76LhEk3pyARhH456y9Xb
s1dRHqLjDamlbEu3Uvv5eQc2In7SgrmGjBizCS+iwArMrvTuioxsiggAJ7NmU3G67aQr5phUkJ7a
LGuLA3QTyH9giCVKZgSMIlVxryGATYxA1i5qYwjccuby2MKLWFQZ/gUgza+1S5msMyqOnziLj81h
1CGEL0MS6SMZ9sWHq8E5XyE4KJvuo8DF9BHxCnvlD1na9/t5XQLOKoJXprYmCtM/HvGii/Us6yVe
ukFiiXXtv/GUCSZqzFX9SN7OSFaafHSNNTMTT2fW9ojnso/HcaydRbz++Fsj/2+2lBhMuyAQhV5E
KgU8873Pz3xIjC0b//CAxJ0r79VD7qzphb2pLaJemqiIAtTBU2HFwux8JdD8H0YyWHLbdE/h93ZS
BCSuZNAJvw+KXenfqZ3xLvNkmN+8cPhCpEHj1SauUG5QZiudU3vd0xTCoQzc89ND4yommWZbG/dF
N6fWfCQcnE4AP0jigjPV3IohkmC7jOXEIUOWqUhsNssadWC76vQke4tpDPbtUfQmdRRIG7uBTHlk
1o1Isp5EXUwVcqw5hcdxB99t1tFRNIA8lVYrJlETe8VSK8kiIDjl7EO6y+dg+hrig/vVRuJ8pvcq
pWloOPWfI9TDNlPhsp4AZHn3AyplMh15kgG/+8I353n/tPr4wk4ml8+bTmN83G7rvJToQIfa8SQO
DGhoMlqg4BqA5A2lHOM2f3WPUqiUMBKxAiWivukq9u7zrxatbbYhHIkzmGLR1vkwssp+r37O0ejX
Oh1SeI0QBSIQkz/gJgTPiiKVvno3q0DnCJm9VKnGtBb28k83HKnk66tRnddIU7Hgxryf1Ncrw0I/
olXa/Yxn9ccCdXgJdar6mVLcSA9JW2y2nBw1YHJEOH6afz8vd9tdd9VjSB6h+Gkd3CNXdTBN5wM0
TX0+NkOHL8mj0mQA1Mbq2HEh98lxJP9iwqSCY863yHwfPMUNU9bc3rxtvg5lUbvXwYTss4DU8vZX
C5fOLdC2/KB82/bMJ7n0C7HCFc327l6HtOrNQykFagNcQ1p01VNZP9QBFUz4lpRQh5spVGU+exNu
QIuaeRBOPJjup594wL5XTxrgBflNu44JTtDc/PJ05QyO32RLrrlKmwke4pCF/Em211v4kI0BDe7P
ne4WpzFM9dMeyS4SJrpZYVb79BLWFAZTpZNiRnuDPRZyBHU2729jXgenwpYuQLWIAAb6nrvaGo3k
xPVLdrsLHVYwhVqwQVeob+O83EQzyaFobyMGZQzasdT3Lgn7dU6fPP3b76tj+pte8ZFH1u03c/e7
x3Xl68/EC5R6VVoKB3SQSzXhEuHxYIrUnV6GwPcGiLCs3RuzwoFlzP5KOqCB91MLxGiIlSmy3TQm
5jhqDcqEqTPSriI4bSzIetMOufPW4jSaYDZQvjCVzheV3FuYfy/J1b6a/rpuHBh8VryOfF1AaF0A
LhPHFfdIIhmnL6bVEtHHvxo71eeV6CNIgLT3sY1LVdptZ/6DRuUyAIZdp7N7v0j6h/HyPU/uRzBf
57Fa4mDQ0AaE7DBgMDT8XA9tuXSKgKOfg5yEJQ4yUoIyllRwbd8Xj/vzmOC6Y0+M8GH1yttjVfwp
TjBQvJa7ZEvRbLWR+FlodzuYhkUxDZypZclLhpB2ekUhmTR0dqscMUIe1CJLa5kfO32eK+oeWNYy
zbNkn24oSvwvHh/30WC256ggrOi4sMM0aZYcfN4P2ggGwe9G2giIDGdE5MKXT83TRud6JBEua5ex
jKS/eOZeoSvaPyP1VBeaxNMHs+9YuNwiJDFMqjLWGc+gquzHhTzB4vIy9o3JsqjWW7eX5MXcrU7j
USMrhP8h+qCP4zQo87m3cxghj7v8h6lXjvTWZwtI0sROrw81/BJYqahSa6B0KyMIc9pQ/EMFEzuZ
7kW8f+06wV5MlY7Hj0i/9jmdYyabRzZyfDM9KoPiwIWNciXmv2pTvNDbQ2sO9S34fl4s9MdkVbVC
Q8NuNW+vXGnfuYtRqS97+7UPsvJ7SEzaQ2tYWgNdqUa86f6+iQ6buBrH32dfzaYlRDgU/lc3FpLg
8WVgYA6cNf81jLTlhWTu56u6+H5Bn8N8FXMnOa09XPuke0MqZvDP3Kzn+b8v0jVH0hjSPanpINvf
Fi3deww3hmS6C86zICm7QsM2p/TnoZdldOXO9u663BE4KuzN9DmV9KpLSWVR33VFEkPO8I0MyYk1
yhAFqJWx5yyN7zdHnuHcvsjNp3JIVTm+AUBYlIDFM9qfvnAimjJ5Re9MJ+1sxSWNoGyc5R7AqsML
lxBgPC8FcaTOynqdjtSnPxlJNV6apW8UqhS5LKXvJEIxvj5WX24+wFV12fdWy0oaMtte5shRP7f8
oU0kBiqLaEYpf9dwHpR3iLHBoTz39vxOrIxDbc4yjRyESTrkHUzkyrYJvaU0tyBR8kN630O3Udvs
si224uKE4rED71fWRLy0ed2Dl9H22Kb18j9Zm9i7V+aiJCPppr9wl9GNvxyX4jeValTDZbDqtSRP
fottSlqiVsQWsr/luqeqqkmSwCanxMpWlvAsKOQeclkdC3E2I8LOq1WWsWjbmN1aPNg+D8/WWCLV
Qkoq2unBRf9e/2DyiqqMKTvT6vtZEeeXfZmu25vPu5LAgpnSq4HzZThpQ1VKEhUZAc6lGerAZeS5
4Y5F3nC4ig8j3j/aBVfbS9ymqe4lvvN1fAHaTMI1XokuFIPT/pQzd9JIfqjOeLTMwAdHyCn8ZfCu
xTWtZtw6EahDJTOraIe1tT4Qz9qnnLrF/RCyYNYEhcBKdambJeEiqyUipqqTIpOcZP580uafVxls
HsHDmLkFamffcdQrwxPuOIC30aLl49XOG8LUtY4dw9UTwdV6a19fdVLYu4ApTDQikY9s7iRVPKmK
Pkwd1HXn/JxZk/+1PEAGFDyuBwSSSMWwVvNbme+h4x5Fbm7V99uclbt1JdkocJm4Dp0SUv8bd5wD
m6ML+BnQKlJMwv5C9jUfLwFFoKC2Ny6CJIBYp9TOdVZTX4MoxXYZ0jSeJQeUyGKSgn+RXRgQJVJQ
T1fVx7MNVqTMZiwokTXZT1yjyqv8ZDtcWC6wINLOVtrixg0w4kEwfvzeGYqwONvzptINj/jQNqwo
MIaNks4nzEi9zla4mi2xvrXuVew9NwzjFu2y+Yy/qvi4ep4/8fzkB6suwOAyJPmkQRzZfaTior6Z
X20hGurXRWEjcLM64zBqq0hd4rZQkxGP+/VGGy0Wlf9DRmV+LkWSEJ4sFXhJj5kUJlKnEs039RZK
ntgiKPgBUa8sK+IIBIcR8fA3nAlKUrztZk4LmpK7UHj7vQIYHgxJ6yJhHgoDP9+20VZE9pZWWZfU
5jc7eBwMeE/2uA6HYE0+3B67HmauMxmR6cRuYx9hzGm57GyiRoj4gxRl3NG1tfMNzpU6bN37qisM
bbX6eTpa8is5iOeF47NHOXyaEcN5vCfCG+XBnG/Z8uCQTrgbsh+y+7uqj51uT/65twDuhRvPFW1X
uZGEvi1HAY1lwtg6gg8zmDJzhphh6zqLdYdhiSS6nuD+ZndJAu8hsHqpk7feLO9YnUg9q+1gRucQ
HBcNUkCmzmFEIx04+LfI8nn3mxpitZbnCeBnfZH5/BdQLBGQuH2bt8T8uAh2OxytuxriRrhF7GG1
wT4TRZFzJyrRp/nEMJLiBXH+InkE8wfZZV1a2LwkG5wm7q12hG2veD9X7/MsGHHVaJAaV9HXjtvr
AqK8bxj+mavfP9FsxrQhU6qb7KSkf2GjXy/ZWGaM8NKQv5WxuU1foEAYgiiL3NkwNLR/YmE20wlU
ZtC2kQGWbPLUrDGF/ULBHrrO3HPSk/9zZrQwAnp4Ov/OfJCjdLoV99B8eC1klrt+eflTEOZrSA1c
u5DAUc93eRXbYa9+DNIpbyUa+pgyUKASGYz1tLBjdjSeJ/wAd2PKbQAL0ssDGF1RhLgQNBi8748p
WGgUwws8kPYLZJmRJLcQTMUYaWPurjccfsuu28zTiVebW0mlpc+xUQyyNtW/FGWA0gtSpnocmoHI
hA1bcVRdyuap10w7J23p+I3Tq95NGrvrniSkaNhlmQFkSo25l9aHcqPhVnAwv8O80bUsNeCDWDR2
Jub5j+G3JZkaJUkR2dEGKfQhzlo0hmfOogPnIAhrZSFBJnl7Ju8l4ESXDF8bkRVYgreKxHX25xu1
B/4819yliz9FSN8nzSU1fnRvnpvAkuXp031sU3dnNmVHUPhtURhbFKGTIByAzSwZPwwEE8ycjpg9
iXm8RgvbQSEbq/Xin5Y4spFDKI9luJScoapBGMSBxnKnbsWHiygSp+gyE6YFy1LkMIkMVPEs8pxb
92xKskD3Rzotxf0O21FhzKpWHoKzhbj7z6OlKz56tKlaBBNnxB/mXEhZlaqmjTGBn+E4W3aypRD+
8/u+xbtGgUYf8rWzR71JOJ5SWe4kuqFkbAsGPsUjqYRY1OkYtO+ZAG3eO4bjKx9irmzRxzftQECH
sXsd/dQi8+OqXy77FjBbJwsUe3KdfBbz11Z2bMwkcbXCTTR8x84Muq7/uKYoMVXj/xoZQ/Hw5aal
K6Ht+8ZMKBqU2tIpdwwvLF2ctGVP6lCeitipj6omchJyfNj1z/n+/MXBxdTiLiLZ2pN6ckWZJ65h
7zHUlyd3/rY5seB0mlSNkeC7fzQAmoe5D2Q7hYITal0A283UBCHFprY31KKtHToBrEMlRmdWG0Pb
YlCdt0lYMBz6NGd/hJL/iWKsmUR1z3gjPwUahKHYeKl9LJtD8qwXCeYJM2z+4iw4EmvYYDNPuWGD
PQThhYzA2Kllw+gGwcC81BlxngDyK4vpzjCTUZbqZBN86PDNFRNtotO1eYU4dJcQpZxHLOHw8zAA
DHbTK55e4+r+KopfkeCyURjXVb5LIv4YHhlfBr6QELEGSKW8d3BTRU+QONM+KOl3X9fd2rMDTdQd
8DCF2X2xCfgc4HiV5KOjmwT+/ksCePUceQ47NFa35AXi6EbRPsWktjSyVlvugcjwltShg4Uf/IDR
IqAq5fAILlHrts/PSjknkR1UpjqtuqLBCBMCVj9kwEqY4VPSdsozjsynY2Ciyeg0mxDiJh4jHsBt
DOL0NrcVRWsyrEz2hWw9NJcuI9bGHWYbBTZQ9O/i7jYcYH1BAue6ZxWedSaR1oSn/GEfgNzSU9a6
PKGIpkTyNVOy3RjuRgzdfALYg20hS3IaaX2IVXiI0MpgvISFj9o8ZNooIF7u1prVkqKlZ7UhtLnT
e5Fj8inPyWR7NyJitwDC/KvPiFxOorMqXi/0B5j1oNlMYBjPq6DEb1oeEFOGmMsXR509wpG0ChWf
/dN3d7FZfTzFQ3Fi1ZZzcpzNSY0XeeE1iKGxH5ax1+MmPS72Vm3hFkyxOVM7Pzyjeygtu3Glb09e
Di9YgSpexwPu3ZzgYvm/ydV5Rac5Km7LN3hDET6B2451IezbOm1gxqdTcBC6zwgxqyRQp/22EK6F
NKSGNb4i4fm3NYtlnQnG3Zri4h4gCx/rdVIu0FZkPBtfKd/6ikbVNN5FBdQB0aYkmjWSfwDMpI3Z
tJQjJx4MrGuxZtuBt5ptTvd+fhPO7fh+bO/xatkvdBrovNOcWhYEzRbELGwtLL/4EnjazqgTO5j1
MVlz9+6qLtdeNP2FOs1zwD5f5IdElfCp7Z4tAmh2lUVsCxSxn+PsPZFiJG4KKD0QjzzzgxO2WX5J
9K64+icBdB9sGf4VsgwhFjjGBzstE72KzXPNyrvMfoCw7k30WVkWzDOb0XE2NY0xeTlWHyfW48PM
fr3r7ztgLm7mdGeS/W3mC6HL1LAHWZOeU6lnOlcdv8XU/1+qhTVdxjj4c/v9p4Nov+w9wMrFU+dP
tCGBTjNOHQvZVftx3lmJLGUGrdbmDIptYxIZeqIGR1sgiyMoFwSIGg59s/6Hs4ZDiG2+GI2KBKN2
eq2rbdcC3e+NZpngOQh2alsWskhw8JlCgnLdfgyioF2YY5toDTeDo64fIIqm5Jl6iE7QYb98WwVI
R0w0zJAOzNqyzSuLQGPAE1mWLEfbkDxxqQYsSTnoWZ9BH8KeXlsRtJyjJbdSJicvRHHoRShjPj0M
j621JlmmhS8YCdy3ETwKng+LLyHcNq0sY/v/UpWrBgxiSRqFHXMwJAUvgqc9UAAqJiMb4XW25kIo
/lqtuc/D46IECePtttqA29pzg9eeUFh/0rH8wNFoMMzj+FLQlz663yF6fyXWHOFG47knE9zq3lah
1IIJunI0z9DzLgQHDTXKPvgaBL8UndJv5rkyjJ2JQJv5Rvx5Lcf2hl8rjS0vaoIjzCLsUaCLtoov
IpbNmhDNpVp5tJ2qkQm0Wq4foC9C3yfB/dEu+a/CLbhs6858XQmUP+Id9ASgmoXaiSphPRZBXKEq
iZXnCrsHfKlhaQpN1MdxFyANJcgFVQsZ2nI1QHmOLQMaU94ZbIIq61xXRErTCMGecWk3+/ht5yQM
73ACSqxDgFF2/8fhTLPbCcE57fQd8qDoBgBJZsABIhJc1UFnJeggP2moGMXBA/74Ib7C/4TjD4d+
9cNVioRrjZ3dHzGpTwTmihw4/Nc4GIkCvFkSsvsmXQsP3pkwBIzCAKcDz/mvSpWaWHkYobJeDTEE
mlzNLUmevjPP3R68CGu71XF1lr/VhoBJ4kcd3F1EmS9ettXomdiSYDqoQWbTpA8HPqLoMyFOb7P/
WfD5SAJW8FgEZKMmpiPjdckRTxZKRvoYuUPd3mFV/NE2uEDCnBBkPFJqdtc38tyjQmueYBSlY6OZ
vaETsdbdC0rWw/gEQ+QaDNvRYFWAJxobtSwNkG3iVRGSdpvt0HN/18xpI3WY1jgw0n60GxlkbzfB
HS6U0IcNZvUhfEoGsfFdXInaJ6bWGnKmQ3E2fUHA6h5BcdL+KZ/EQXJpj5GFxwfHBFxHtCURfOh6
RJC6wyRAVFE8g/gTMg5FkCec/gj86yTNt6i0Usw/CAQUPMMzNt8xE64ukVKV7fR2EdQ+5krro4ew
vGbEDrixwKQ04XtCIRbV2dwlymI11ClgD+esZwCCahS2XprC9tQLsSAPLvDPcIqGaAM3s4YJQsfa
fC46e4D8xsx7ZcfvQmfj0tcesNbBYbVIF8mkzSYTQLsTLmWysXTU9CTin+qK/SxFaPLlTbeGdFJJ
28jJC5KE4StxLR5PEfbB0olkit6xISw3JQsTfecN2/pck/VrkSetTWo5wGxK+B+2PXff9xH7LRWm
ZO1fch+Vp+MgjhAbTJR6cDz7B6eF8y1jKZ95ncHBJmswq+pc6GRlX9wDvTq8I1LsOZ+Uc/APB3Pn
2qtF7nW0/9yyV6v4BNzpbaRZcPZYOM4OBftDoFYgk7W6/87aTbeGYq0nd4vcXJXrzyD2T055VG0z
GQP9/6JAMzQUHCTAT5dsooGeeXC+Rs+wvApBbWXo9pP2pCbKE6lFrKyaormhwMrbl0oZs9Yd/1ol
+uflnBwOsz9HuROwMVXEWS3uQqcmHI/r4DJHqdyyGcr+6uzMBUvukAloJollgu4qD7dDD1OA2hJu
3DN1lCBowYHSBLJk/vWncA9p1XRzftLjhdCLaorjqH6WbjWUPUUHev1WbnNjZ3AbJdF7zZUUQJw1
m5fENB/RXqo/aF/s6auGNmEWbpBu6yWpEG0EW1MwCgGHItGxGd514QMLSEcLNguATtd/OXGEgxpZ
f7r5o+roJMNsQETlKFjC1SD9U9tPu/h45b7f00/jPX8YnekuJIMppIAC+/MKDx/7MZlnE517HZbY
imfbBJh8X4MgE9sUBOlKzwt3Sk/q9zvj4Bsogi/gtfbjuR7YRrC8St8TbCEZ0Du/GxTbY089NwLF
QTKCxyqJ0okglO5lw0bH9rTNZmbTAkkFY3h1B2DjkF+PboQ9gWUa4jx2X73z3kTfRnxe3CBVHwKm
DeDZ+GBMDXTsryYRyDeYE7+BC+0SoSSCQGX4DyKlyC6xMWeu5wImTHP4gljU3ZJtapcd96vhQXLZ
fBoA5vCnK/sveC95QvK6MlUXDtyoSLXqM7VY2WebfqwU//iIErE1KQYMM4ZhPOsOgGRP/Lfc0bnD
VqlYvjOJdRNkhH7O12X91k0++kfTlUfyxBBe4TQrnhXbl0V7Slk7fgjFc1HOfWPUqFCIiGf2kLZe
D2ZHvQhAEoVO7PfCMIoT1j6n7IssC6pKh9/Mfrdv13CukKmF6llX5MJKSnbxntYUaWpMSQ8edYbI
CmTQBjslS3pLAWdYPpQFDV/xmidsPURyJaAjDzOEYdlLHs5ZOhSc9K0Jg+iQPruyPBPUKvHF6ldW
+xBpXq1LayGmAFUoFOuYFZeDnplNxzsYZzN64iF/d0U1ac+kRWyoIXf9MIC5RS0nho8qfo5PBDxG
HK/QBE9AgWhTUkbavgYIPvUGsQHSQ9qutt+zeN0OJnPiDbo4NJlQcoEmzQkrnF59KeFv7x5p4V47
mMEpP7dBX6uppJtbfBh3Om8RZsZDijA9qVzj2tmoaz8lW1BA3gv0nq440M9WBl9NPcqztWFzPfCj
3v2W73eCtyR3BHsuRho6atT+XtPrKfChNXMec8zOzGcfF3H9yu4M8ABH8eqqdzx7UBj/4MDd6Kyl
6E+XSov5VDMJuwywPng73MyI4CK9IUCPgD1t3Z+RDdfNMUNN7aPU0ButHZbSEHY/M64bPlbgXL73
1GiUQSCitt6TAlBePZHIC7a7O4hu22BOav8QeEwA2+4+VfVbW2tTYWiBngh5DInoUQTUDoUnUdMi
cqajm7iKDrYtonSVZpMkgPLqxgozrfre7Zrg6C8JFFOvB6qOgSQtN6Gf7+rfFboPfOVF/ytAl5Oq
4TT9lvUFX7aSyjfNDVDs0XJ/hjmcMBJouJ79vRGSQ4EBGzFgQ6BQQBGIGIHEEk41WGETjLHHuvlh
iOCt5E2VGxBdfGpO+dVO1N/zDvKINeGsrXTiMoCkv7C9ut5R/JFe/TDGXmsSkSIzSCkHpMqu2/pm
BJiXbR4RPXwrwyl38py6kdZQFqTxBRvlTgrcrP+eLWtxfWG/HtxfZEgyIg0kmf3ALpxfDE0F/PcE
0Cz7ym+fpL12dPudqMXMPf35hNt+y6YK+i0UEriceqWU5SOa4n7HyaGS7Lu7s2Kh7Ev5IIxbe79B
sw2KDn7jkXYkepwCpSeAEvOxD94vV04L7KRbp1m4Tqas00kSY7NlwczPTIwGBdm8Y4PyuwbMO6G/
ODz0DSquL5kHdB5Q53HMeQptS0uzu5f2y+ie4c4JpU2uJIhxiHqtQciQUmukNM1VC1Iayj0vuKH6
6Z3AAtivI80mHol8FAPqD3kuWyGe0LDp1V64uYVsXy7kV+uH/8/y991Qrb4X8q4xV4lSG82Y9GuG
s3z3fF/3oRQcpIQd87ndy07SivN/5ZAALAWylaUl0Z+dNuiPkwJWjNvcUfy2FVB0bPPNlaWhIBgU
Qs6o6uVX1tNnZvh5uIxn2fEkzh9YfxZYKjQAHrVrfrv2VpmOAj+YibVOFVsoi5EyIYxl/l7ExRU8
zXngWX+2XYMdADDt13uXAZrV9W0fkM0JzUNRhaf+rNblA5Q/QnC5B7QWQdlHinPuJSwTG9um3vNu
5aDOdF7oQXD18m4HVhWVjgN+tKtwdWVnmjDUAVggRK923UzbTYhNFI4n03tZ3IbR2diQYTzI7ACv
pBFTPsVFkotRaf6P8YCNinMtn39ctAlopp60hGDDFVWkGr3wLv1n2pZUfz24v7epojpzPNAhubHY
LvWK1/4TUzrKfMHTNhol3opvXXevJWeD4J511/G16PGPiJzAkTtCZsqPIYYMDVCZPJ2eHRIKUfpK
SLA+KHiFwBOv4H93nb00JwZX3dImO64Rc4oqYJDtQNJJlTcChK/beGQLRKvzobnK67yWg5+PDnVj
r3/SZw6Eix7jueBpu3St1Ul4Zqk+XERKJG9Z0BeAIX0j3xY7u0M1plAaPE+GVp/gC4n8T/d8apYg
7oA8ba9ww4r2enOR0ObfF3dZDj2MMTCSsMKPFvnyJaq8SIcOboaoqcDtI9yFBBjf8J2C8jMUhmiB
FiNEytISWknQsntb4p2A+h4DGaBR1TNB3e4nci810SDPLOUkrDxydRLqTnDqAhmT9zGfcaoM8meE
q97Rzla289+ZxPF5Exf0uXmbOJlzDGxuVYk2JNBddmHAsybPBwTCMhobIx4+kCp3+kVSoekuEsrm
v5dhz6VMad+pj5hCF1yqDHA/chp1nATfMrAClcX+AZ1hfzIFFMj1FWBM4ZqZ54UaqB4xga/kF1CI
KUtwCDFS3HkbATcKPaljaHJrHwOU2hAbmB6ubVKpzyPAcY0MtMRfO3dySVBtrFql0oi61oqioYSC
7weNvi75IdLECxEP+J75ANkyje8/KOCVH32Pzwg1bmYgmvno5zUmBGCZA6XVWyfewJcR6nZYW8sg
LIl9B2RayudRnM22ZAWpsZeRAZf6aBOw7Ml1MFqOlUYhL+nJ/idEx6nxwbNiDF/ipwKI/Shl2Ze6
GYAhXD27l9prpXXVbOwvo/8v7hLoHxSVCUg5XTiJ+2AYGq5FXYh72rs9GcoFC/65CV0F1rj1dbul
7E2HtcolM03W68ajoDxQ4YHMreXHl/uyPM/AkBOHSgngmIoSRNmvXuglo2qjB1u1P1YLZ2Gugc5P
sLgeyGkAij0aNSTHAgcBh3FAFHhMOJOUDZ/fkGvIpco7/j6eVj8hy2FWW/IyyqKk1gmIh9/TYfJ0
kFt7mioydSdW0zQpdMxaurZBrFYFcSaoNXFqiTwMi9WWplfeh1yb1nHN0Fc/1M3LHMvzxPceNiCQ
u7Z1jgxJcZZQLMWkrTog9/y6jAR9MmSAk7sx1Z6upzjbSfPia9k5Hll+1MOEKHXS40H8wieIul52
vzIdzbXmUJ5y9WiIcsHmO8Bz422wqghHpdGpsHZUMgirQTOV4CPPzgp8ZF6adeozy4A01cjNSJuI
HwwIjE+zxJWp17FUK5jnPRZh3GoI2LCOFdfl5URmeCp8hU21XxmuvXPqkFxcyFpVDEpDVT1ge6oI
q1Hx9V1AnzioxIHZBPx6atugv9tZ1qmeGmes3KVzEyHY7oixb7PHTSRissqIRbtquU5E4+G3eNKs
lVuEzGu/nXITh2wtv251+9e25zeLRcJ3Z0wwXZQU5eJwWS9IpLPVNMqVgQmZjc/fx5CE0vJL/eJP
+M8wBAupcSI1Z0aCLzx8wc7KVkAPVxTkcdwUnu1hbi5fFVdnhYkDSir3ulWITbEeUw1N2mauoJYF
T4/TOcl/7Kvy4yA/S6yjr+RviqP5yNeUOBBdG0PqQjpeaIF+AqxYgIClf6xF/vh2IXq6EmSkTsOU
f3QosdARoQzhFLuuMVYGHG4mWgvGL7E14kibOTNwpVtr9NLrMPmWEXK+XAphs0mHVafl80Lrvw6B
M1WoLJl/yBghX3gigK54xdcjLPyNDflNP1za2sfummIt/LvrPUuGh/GW6nQRLNcd0wJUahe4SS2e
j2KHVsMXe7gYJMJTQ5+vODGZaF9XcR81SLjAyA6RDlUkTKzKK+KKROZbkW05csOArSKYe/OitY8a
L3+Achngl4pVqsb5wFriPLRVrFZj7KlA6MK3ansxOe5M6u8zk8wRPVc/zHzqLZ/sH5puFg0nURjY
pz4Y9nhmTrw5IRSQgwEGFDEw7jCNcKRChxj/5jvNcRnpYXZKmxIHrCF4ZaMvRY8F2OV+cHiM8GrQ
1w4ccTKcabOojzpNYDZcoWykJuvpaQt41iTxGSfq/3FyGnW/xTRUm9BZf17dCPWg+inS6sEGlmLQ
IFBCCcwyjswb4OFlMtKRYUPPPA7G5tN7yILkUDsiXjndY7NEChzmZyGAgKKVCvc4KFMqJvJe+70K
NKRCpzFH3RyAUBsCZIZ8OSlJHTg/YfgZ5IOYWrWOJDAsVExsIkyGbxrtHjdFkwqtE3kMq7PsTIeh
rz6YxIGiMkixBVqlfok59c1dknaR5UD2yHvtUae8jUgUpfZ1nG9XDaLhTbsU/GfpGyhOAVnMQQzo
3fL+2dIyMzHeoBbyGY9XEVvX9D4uDhhOwX3rEJ/P02rdhnKe1BsoWC1Xj0K9RNguCk9SWy0hIf+s
kBGRZKFxmL1Tjm0eXYNFWy/orihSdEmZKxTXhOMtekg0DOsu0sEcFxcSo5bNXwk8xUA2RWfo7+jk
nvbyoo5DKo4bWuDyqCKVmm5D9w7AM775GSUsXazUKFn5Q9lu4io2G7AQHzOmJBwDKOxuZmP8ekMj
3cnBu/a3X88QNvu2ewJfagwZQeTRp2NgL+q6dFTGXnIK0MPmw3NjSU5bnQ2JHHbztlnfo8Rj1Xjh
b682WN7Qyc1izL9VP5yewKtNXKCNKO9EHjINzN3sx/Y82kuFDWyQqG6SyK4lAYEfr6W6B0onwVGY
EpQgOEWHG8sJci28231n42F2w0LaiEz8eS6EnYJz3qS1OgqFjtBEdKfQtMTA1AW1giESFeotRlNu
XON6zTlB5mdZ7w5/2mlKg7lnJRKy1evX5Q1457/YOgIBks+nLYJQ/laVQHlEokeo73JE+oo656ml
dYlw0e/WlI+LVtoN2vDlhNq/DtERjzR4NKsGo0dU8rAy4RPuAaUQ8yOg+HyKf5DUbPH5TN4Z04Ou
JgHWfVta2L+oUi3rWRf0vLuvqOlEnbT+6NcWV9zbIzJlJL6ffk/2nYm758ziMu7SUQcRtCZ3tu7B
uuAKPBWoObK6PrexX/32AUkDXfMQVTCE7vUu2UU0pQJlmviZQZ4XmBUTC0BTEWcS0CPWHcPG/wTB
yew0cqCoQ2R5q1N9lc+fuKWLCF5c/UJU+KOnhJ1T9MiNYtHbDQPRznaSm7gyG5pmjfvXQahi4W/k
IRNzeFuXqcJvjSRrSGuNDbmQkiJUesIwe8ldnWJQEagXgeAmhEIUNmFIBIF0/WKd59QyWbvO+OTk
3lT2iysO28ptKhOUbnwEGiev2hzJu1t5RF7DFPauw06PwCrpStulhJwB4ghA+Tb/XeDcxjvPyKzS
u5rSptconVzP2Fjv+AqWSQnv753k7UrKRlFd6HnC6IKZ8iiaHfxkcrnsW+XnLMDLiYqVxiAcOo4c
u9BwAVO+jWrtq4Z799taqITvAxPbc2Z8Zf3b+7PeJJPL2+iGk6Hd3zkHHFhSPN4w3wvtJuiaAMnH
afGsuK5sEiH/C1l6iTpDEkj7CeAxQ2M0HU2GdY8/T8PX9LNbXCFRvUhdevOYaiOsFkV0usEYI/KD
JZi4sLCFOYfUJ9gyD0DxuRgB/LHH8MLDegKvc6JckSabugpmf2OBwby4GrjVtH+QtGfc81ISkiIm
n5jYw6hfl4DTzNy+7vjhkFYQHokixcJ+ay1vaGIhSD+qrK+b8KAWkdKETMTgCFOrpQ8keNe6XlmS
HKvPherPOafm65tUxGkzkQNEsFYJFigAjuvDoXw9VIeH0BW69NzPzN2n4rKSXqvfOQZECgj/TbNg
PoOPp7ocKta0+oRq1FFCE7MDaFBOJARCh4cCxbPoNJvw7OiY6HvadeuXvp/gLTAhm2QrGngjd4bF
b3uGA33rYJAbvLbQC39loWm8DQ+3ykcaQy2JJ/QM88Z/ZsCXnrVoCByeG4jeS2NdfSd76Cb7LwGw
4o1h/zGYfUkg7h74g3J1qIi6AFXJhdrZKIuhEi1arf/TG7IqkjTc6BGInKDwXiLQN6UFOIFVGyEP
mdr0BRXtLXRrb5xDbvpmodDUCL14525hGA5y6vmGgYwxRccYi5tJkmb1xp1LOrpWrYVXZdZ1A9fL
Q6EdGlr4vnHujq40PS1JqJ+uWn6Fwnqq13z3Fas0QLvj77j1qmPnaYMUg7JDxIaCF4zagF5hWNOq
C5PybjU5dxK3M3+wMj+3D3WRCTBFrGJ40PBI5Wx+0wfWhrzoHDeZ/O+uUl6AMgxg5vZ9IxGPLSy7
7Qhc3dTlEviNINGAa8ZAP1/AN39BpypJmvVUSGsXZaJOzu04NwRqeBOYapFoqODups6y0jRt/wbC
17lwpoAzJtny1c3SV/6qgbwSGHItHsDtDtj1ltKbLS6NhRNla+XeHMOaEeV6kVDhNF1VHGG8ttZw
4QmRaH83yRKbeUWuU49hl3tbGkMsCVmaWUAnCjskqSJCHv+r9SAvckmDhdFpXxXyqgjLgiG7ianV
vL9yT1WR21NXlS4QEUFTmK/vbnifkfhg6HTTuWykypLuRVb8rhs2q1xNuZCrbmbzk9cAgT/wazF+
gtJpjcoKxg7gvnYPOvrSNhZpbUJzuE6/b9O4shXTFF2QBV4k1dr+CPZdE8Nal/gdXeuPJhEFAMW3
6grdR18+pIxgm9uzoRridaZYqzSnAbsTCbuEy8uUaOgRlLKHcVkVfQFbiHiHQw2HJ4vYphpaKwpO
gbWFD/HT+osIWAVNZNYq1spxe4+36NXUsvu9IbVNSYMwCeKE+cmZcYbFWjW5lJ4GQ/PXui11dKz+
aVQnti9bUz4Msn8+gzkQ4eI559TYsokRNQgV93YMVK7qF7+jGSYK9SqYHWqkQjN30v5A8BTVRoY9
AMUa+2Qo1Cgx3pWKKqaz+5OCdzMRPi59EIxZ6hz5rwUscg3RNlsKWg3aaWHuAOMr7OmmcZah8Qsh
OcbANYA5YPL2oFrSXjpw2bZD+SdUTogRXl4USKIleqVov8upxIT6pGXOiczV+A5DI4giTT3XPKNY
rpC7NKNrPX7wy+ghlluV0RoDFsqbpUGd2IthAXPDj3hu06v7VWlryrqHERWnPr4dTIve0XVyHlwk
iQya3SZzj+XhTslBmHZs0rZqNUWBATcVRkinRxcbqbiKsGhxymf98xnFkTS2cCJwvKZU9oFT+O5L
8/PQte20TMCUvTi50wlQlZ3jSJCl1Ydx2qlAq9teo3RHofMR5v4/PRMv+7cjG7rJ9SvD38cq1k1f
EeZdViUmI6obzXqx1SBtESVw9lhf91X3O7xgpU2zcLui88UPzeqIgNAdshiScctXdMpvnWgLz24g
SAfQQq+E2QLAyswtjg7Whp8jFQ7jiCOa5ztgOp2S6JCndfgHBO2D00OpOlElo++Msuf8tHsUNJYH
3oT1R5Ods+ZWen/BK7tnMOv3rs4e5m7H1+QnVfag0raCGcmtttYPUb1yx1mxUqjGDBbjmsEQABQX
uMAixQlXZ13/wXRbjRnLzIUTda+MNMChA2MYKXb8zIggYJAVMVSn3RpBX4DmbL26Tu/M7liQJOfg
VfqLI11tKwhva8ePEkuL2Wpg8B6XVCKUd7BM/aF9rDu6pLs7oHdi0R80uNlVUf+cjeAwK6EdwvQK
VC5qkDz8Voi8+6Hy0C6UiO8PK8atwbAOCw8T75cJ64gu0n8TOlzgUbCX8ojkOf4kFj99dvhsG+GM
yiQY+YQ3q99sxefw9fNjtfHKGQ/k+euOHW9DzP0K22G0frX9RTWeFePVqZXmj8JWjOpNaR680yTe
ojRIQqSU8K9/FeXHZ/bOWC26F6yoroB4KiJXplqTPAccHu/cH2rDtFKrmthSdtule2tBSOu5jb3a
+DKKHtNeHrBfmeNDhun073o9zx4JkLZaanuUoU2zpuD8aoZCziJC23AGDfqEa16BeBkld8/DpRNl
L0EAaVIqYnc+TOovhrT0IcnFsSYg5MqkKfECM207nGoJU7cFU1+YqMfhUJD0KjmyuC9sy3RuUfYB
JyRdVltUPMAgJGkKgE3CeuzoFJiGy0Py8VDqHNKE38NEHFBpN/N/W+T0xGxTwx3qMKm/k2x9CAtN
N6T4JFOLo2HZtwG/fA/AqbTFTaNjCu+UawXpesLE+e2Vir2SXN/kmQyFydAia1YMbpI0tqfMCLS8
WPsEd+yvb7aK6dbpmhVZBdX2KfeabT1dh5lThuHPamplcbQLgk8xUFTk6ikgxQAENnkXkuO2y9YZ
z9CmI4APJQxllPDUA9S3DCUCrb6a/stoM1++kButprwfRGIEA4fRhxm+5OHBM9Xjr9YZFKcGnByU
VfB8s353i8nLMEf51he1QFrFg8xRXTwGm8l5O8xoC1E00ALPezZ1yfIlTQKj+HghXR9tklPr2OVs
6kjApO2XN3Dyknp1WEYvGek+DlD6auw7QM4atqL4XfToRBeqLTxmUVuA7h+ul+bWIceI2gnhghmM
F9URxCi1Z4vOhfiR2yH2hFrVncaGv2nvEzbUUJQTEoHpe+34ky8qmiwjrX9JqLzl7D7aL9Hbpxp9
kQvQg7VIvjZsrbH9Y7ikoh+ioEvyQ3j9la81M+CqdPnohaVY6kxe252t7ok/zFoV8P+ph8kqcr3l
lVFAGLLHrqUQUYoTcY/WDbxOZKxUU7buZBopynHsMnrJjTHwcpX9V0LMTr5U5fzkTYUGaCTzG7ht
e+ZkhdER6Kkr7XV5+HxSRN1bwjJfdYydZpMxQAY0oCZuInNByuzGl6xLKSbqA36mElKIZK/G+xhb
FVfeG1Wawp7cQposUOcv2Bib6J0+avgAgF1IuF1VJpJmn+TmdFSxGQx3rSYIC88s5/NoQwo5zgOl
Fdz5u9u8g2OaX9GC/NEp4msoL+D5a6Nmv8oAWm9Yr0VU9m2JR3QjeCR86oGD5NMLxI6rM4cyMhMp
B/1EjCaDGiNHIiTYMymmXJwv/GAdW1WOzJ0i8KLRg/Ae/3adcGxiau/QW/z2XcU1p6S/qebqKTuB
4pw5+/7ybBADswPJSeV3ELWqsfDmI623hQyd1jpq5Nog2R79Q3PCbwXLrbRlZm7ZguGvkjBAXL9w
7uR4FQWk2pOcqsrgX3k2zCKH4IS5/Mng8ZsQaVpWkQzrvjcjP5z2GH7uFSWmnT7v/Y95CV9gKakc
3VhSjMaSZOdxqVXz5bKuDQuijYnEHtj3mLjWegO+QyLft4VpJuOYAViUrulJdFH1dpqHhFNBGrz+
iEcFw8ERnP+SFUtE6WBQOagCyTM6VilnB6W8oBjBFuSPp8JOXvrQDjCRZK3OFDAJ4HbTBH8+ifi7
kKvPh4hsLP70eW1WOhyMXHnLkyiCiwkxRwuRDyGBXJtkDO/6kVtcesNeSSwWOphZejPFojC6rosG
BoNoVtVvB2FS2u3ktuMVqrB1jq0KAN9wmlIed+2H7bVpev7Vt2ZYz0Bjxvckie84X2r4UvAdAdvd
UBe+FZUVFvnv0quX4MO1crDg3xtgM+eDIIaU4tbAVWeu34bJCgOC03paIf1u2MTdKGqIz6BSB5A4
h6YzK3u1prIKYsOyTgX6wX4dLffYxVnY9IOdXNsBnQkHwK/RqYEm3kyQ4XWuqFVTOqsHDIwl6jFs
A+5ATWu/VBY+PQgvI2pj6c5xDW03WBZQCGy0/VwwVhfRRF0dSODPBoAxNOAP31BUEsDWWIkifrdR
MgdimoUq7cSN+Gb51MN6690yFxNb+4Tua7AHUMPZbMk03inelaV5RkmuZC0lgcnnnhD31GFd/S/Q
0aVT1kKW5ouyEknRl9tDd3N3unUh5Fo43MvElQN6XJFvrWsDmqTf2Nl5J7n92EwdG2n9r+/NiJYl
PiL4JaUnwnbyhnLAVezCN3CsxHpdbc6Kg32R2tGJCf/C+KKxe3PMg0nYlwODjJIj2iIDwAQ7lZkA
Fy4Ka1MM4teHyWiQDxi4S/x4aO0x8vmjEXACQHw6bq2po7O/mBTuN06vFaiiZKfdgr9mMJ3+xSc8
W8L81EAaS+kVFXXHjtfGPDlEpVBq8t4wX8dAdDrRKzLt9C2ExPrlgd4WoK9KazypUA8XnFrVtmry
8BbOXeEUF/U20Yim7WI82d3Fh1hXA0yrW/r9PG239n2r1p8vdbD8S8ZwttIULantP3YEMWQPCAKj
EmJ55O3B3zXLli0CEeqrSJcHWermFJlN0suQAoaPJ6NZ0FsD5/RXCIxBa64dMBiieLQ8eLkGkwZt
AF2hsJRFSUq0Akq+YAF/M67hbe2F6y6nsxcITZx8s5Atf3jyvssFiV12xP3jsVN1Z2gJ27jGrS/S
66iJYkjIdnssu/IPjPc1pdghNACwNMGAnk2m/osK3qv/YCpkQMtc7w4wFx8p2V2zj0M4vApxMrYK
v6xS7eBqxoqx+6AD+bGwACRGPIXGj2wtUX/GahvBpw8auvZzHFGijbs/CV0ekWSBK4G/FDh/Ltpr
IQyL5FB+nZ/Pg1mzqJdEUnrlN1iCvdxaCEcJrAD54b3//lvdHayuVJjfYd8Jx7rFH3Q/0EQJ6R4V
+mlk1EAvE2tOeEyPIHyxP9tkMmwn3aNtuplwmofvp3v2My//mEBtCgjwzFxu9qxFlSsA1UpIlZFi
eGG8tFI63YtRXPeXxQ7qwX7T5h5jS+/iIVgqOvIog9plkeHlRiTg2VTkazCgWXpoeqOL6UXYUOIJ
Nov/KAJ+aCnn2At9yhJ8WuWaG9W+S+jH5AwJM/D6drrjSrN5qRmcGmfnljVRnFtBYg5Dm6kaVNzG
sivYPMpcudzhSdIS8EkK+Dx9XqjdE0AmxW+O2EozZpL9Jrma8cwoa3OxJVesVGlg1+SEk69ph1w5
lD2VWyE5Wx/aAErLfeGkdE6FMgyo+yUkTcKTENO3HsLMEazFgMw8DMbPBoO1CcCMKTVGEGxX3hoA
eFzzop8U6mtjyVYcqsedA3GpHmFk64kn6xWHvs9xaVSxTC6X+mMMLxldgH+BozNIaKIfV4yuHgkt
cqTTlGO/H+m5OhT+sw5sm3uvHmEabWw97OLm8p/T4SbmZKs9eXl+WuL/Wndk4L8Wzw/ponaPf63v
Nte/L7h2l2HfnAkAFVWVeLLDEsp0xT3qBB4TkLxU7LSfuSt2bWcpldgzGjwtRFvmYIdew0Jyy88E
ivAReqTJFLiOBsZKT4+j4Ga3/LwBtv4kmUwcVvwBJOPC7FGh6MDGTsFEwLJHjGg18jsvIOCvlGSA
CAhQv4Pns7t8aPaXU/WRrmiIycDtv/vHlBVO13wPaf9PChjboO/+tsqamLOlAqRkWLcGhl2iDDBW
4gcSiNGVz84rQHGwsXtBgz/wOG6kk1aupHi4mM/h+ozk4LxDQP8oULMycRBSLGsv53IR/VcdkZU7
gxwIfPZTKU+0KDmkFuTeY8KNm62Vc9ucMiRtiWWn3foYpJIjNYHb91pbRVvT9VwPWkhggmqMe8VQ
zRwD9HAdTlbjaGMu/XalD7SMH2e2mKY5K+bj2qa2BZvgbqeIz0LHgFe1O0vYbGJow8xSk6pmtJwV
w6dUx4LyOi0U/+ql+oNrjI34QlwR5oXDCNfJr31teZW/1SHeAlzGCP1D4Rdgw9dW0BqQorrRJGNM
lAasyiXcW9jx1CjKfx3W5EETVFyVPoENwepraqZ9mLKW+0sW+3cEK6/0aAkeOVrMjcBgnVCAzjIi
d59Cglbbmz8vZbS0Hn8iMNZ+ub0ngq6aLSy6AlfjRUk8/OSquLknYWYFtGpk8ytoZQJsFBvbvcKE
BcPmEvUoX4y909r6WJ28N29jMxEXu2iBdlBd67PJWD6zMCRM2HTjDcDCdnhFIiwORiMX+wRik81Q
A7XLLXG1vku6BGfrhbozKrKtfLR/iv2CcSHibNaVOep2lDcZ59BHCEtmbvOPOpntY3hCi/leJ5+L
lUCNdn/J67tHFkuwpV3nLA2JrUGvjlP+BYGa7s8PGrfbPw3nAl14A+205t6KOsScly7ckoZ1LrKF
QBaSpu+NWSwqnMEmhgLoAfhwH+3UmFcwe2A9EGp7o8Hk74LzoEnEAQ7btiZZEdCihrSLr6JghKK2
yYOVnCQImrDtJQNoU18p0fRVFn6m1m+9GlpG9t49Bnzaw+hCTu7XkWC6cstnk13TJH+WHmOpBFqA
OShm0CAbpZMGNJUpjrwGdYCU/zIwfLxfxOh19WOOAsgSdwWDc/EA+1lQyfbhA1H9CGXjf9MhrbfJ
y/4NJu8O0HL+PNNFz1fhAb6Vwv2tLg3QiVX6k5ET6byS10TzxVIFAcuJhweSUXWgaATPLyMpe3dY
MA8sPO9bYcqoM5QKnkGy2b/enEV1lZO2mBxFGbG2I0wjbqd/noIJSdt+aIaEnOtUtjOX5zEiFR9q
urZIv+laBmDjhpdqTPttEYvkfCuOeq3xLEzUxmdwFkNYZBxXJs2nhhdX1bEV/ClggGFFLnrOjXYJ
a2Fu3Ip3Uf4xfYxD7hYZ1mjdCMgZ0MYHX/C3z0RS+/LVIzKMQoHqLm2beVLpTR1rtvpBkoym2UKg
LBB3KJlLMkMQFQIg/iS02KZq8SQIHPPKkIe69AsLN7X7s5wS7QktZ8ke7h8/a/bu98ZLghXubNHq
iOqq2JRgKCAxW6QbDvlENoi+VVZ8sVhCE73k6yFyc3uj+zHqLqJ2xKgckfinqCaqmsW0BpOzrUgG
UijFtKmUeCeNuXkTtNGfUPvvvYZ0ZfbH56XFr+hmZympCWJSyYVnf6nwRwPSPavu8Ikbc60H/Wr7
3JypghruY5Vsc20bPwSYzCjKI9lSyYRV5lOciq9NZ5Nx/g1Q3y5bKXK+F6p6n6DVa7w7jcvVoQLl
OH9+P6cJ7bR0NmZGKvo0OU59pN8yzGAVwhTAEiduZPKVPL2XdATsDAof6D5gc/jo3wf3D9uwizzz
+YN3KgWSZxXIg4erP0on4GWZ3czWfkCPJkCEXjFMQSzqgrZYlmDDYw3B2PBcbaoZEwDL+Zj6PpF4
Y/7UOForcekjVsVikg5sqirtsGoAu3wZNc+eJYzx51/a72e4koQjXgnn+Fy/JnEWm+Oga1b2qW+7
YFF4UY2phCfy8e+j5hgAprT4qVgQNvu7VAqbNoR55Voo9RHllbJYBivZG96cveeF/z7gj/DVfgcQ
p+hFZR2qeNh44W7euJ+ArRdGk9GxjkWq/wdr7deWqlV0/469js09PAG2e0/prqSwpKAfUy6TqnNW
3mh9BNdG4JK7WSHEdV3GO7vY/rvaWPjkbIKOWYX1wg/rlUXQUErevUSACYcXApWd1MwldE275r8d
Nv9uSSW+gCyvF7g/A0jgEIycNApnWLQVBfQ92ErVU/hKNZAPkbC2O3otazppSycQR4UimF4pNxqL
6pr9dGzuWdVegoXKJvtQHbwt+Jf+HorR4FyXwspCL71nZou2L+vYiCK0GNlY2jmVjSSPkLVTCFrh
eOUFCi7konWzcAcGO2PVa92rJYx8G/dx3Hk1zaBTz0QTjbdYpmZt6bqg1dq/Jse2LgzmeV52BgAj
/TNLcDwGcFESLPPMCI9irUhUxBxTS9KzvrsK6t1E92hZW2YsmUn2r0dzxO81bWho+RJbXyen7WZ9
xKJlgj+GhD8GUyKuDeG0pFlAAaQa8umCzt4wsWIGbSDlt66Krb76UE8yB5aH7LgQj3Lhiw496phG
mkqV19hPzAFTBWL/jbzAIqYZn4M2c3Ssig7GcdiQZNHtKcq4Ts7kd7sW5LqwQkHywHQ5H4dA4TES
+8qXRHj2TyBQdsCusOzgfdR433u0CB6tiWO/l/xV5LLhNn1zJX2X+OKiJmQ73AHPBB2Q37cfxodx
Ck1UL1MzT4mg0gpMimyZ8GmsHwbYHf0j8aMCVtH2qw86TqKU0r3o+nh6FZrKpDipeWNaCZv1xxO5
cw1BzBWhXABDrhb8EkhcO0MhEouvc12b7NrJaLcG75cTgLzPIr/uGfvHOKB3DyCNP/ULyVVckQak
eCOKu/LnaKI5B6PW/BGb7dau1WCznXwSPiwE9A0L0nHHIdmUCVCT1dkvAbiOUu1uaZHVHnmGmnuI
rNNYbSC/ecMbZzHWYokj3IVnmtFglZP90CgeKUXuOYG+OKZ3fzlNkZWQaTst8UXvHUf60TEic2pq
9S9v9dGrOmdzSMs1Rf/H7YG350fvg1JVmHBtwRG22j+kgw/nD6eu2V12ASwD77qtn48j+JqRMU4w
rtMYuOTrTVWt7KdXPfyLe2dSylHWu0m4drCXR32qNHxOyV1E01d0eyL971deSX1j41mYPAVIzm7S
TcTgdK2Rel7GwHk86Vj+ae09/E3s/aviVCN1UavU/Db83zspZ+HCPZXS+mdKlE+QQXe/96FAmRYj
7dljVyaOiLBsFCDyEWxgqapL9OXlTkiW27zWUtC+ffbAT1OVj4UG8hUuVRvhzuxNWnv35opFlBQd
XuhbHORZfTwVvQhM3ZQiiA90r4IouhNz7oIHvyMmk3inQnYNXrJtH6opiY7/GFiCvMnZiuYtbZur
N1IUKYLZhuryfK6L5bRDYp2FglTmYElJA4WjYlNeseOOPYvrQk3dUO/CeEPqZGvNPBS5tKoQ/Ec/
o6xqDTU5fmTN12mcZaTo2uj9eWOdSVK2Hj6kAQcodKYoDguA+ZDQhtef4WGx61Og0VFty1EnjW5U
H4VuidTPyclcdKvk65+DJv/+tCAwrpnio/0/8ZiXasTC133tFUMgIa11tQ2m1K0LhGrJT7KgERUC
E1YTEJZRSKCec6UBnoCzK2IGPnmCnxS9bNNs/uPHFjngzE9t0BYkNG+w6n5UNpaYRhUfXojnLg3+
t4tPF9Qx5uZ0tu9U7oYuQLK6WItRF9JXWWUK53Kw4cohZWjrlllNunHC5VUUWPm3yyLUkZDo7b4B
QxM5i5mcdLe+URLeNKDpRWeqv6Nt010puKKRu7zw0NiKTShaBkNuYGWKsvMT3kWagDfjQgMwhl3Y
hEAORi4HiR372+HUVuj+WxEyCoWtVIdXLEXlyJa+wHGuu9DQ4oztERCbGPU8frG06rTcmnicGPqV
mZLLFE8/WqiqnqIXE13BbPdgP+F3enAgBpCJaWfcxQ6xQXzCgkNp1iLLgEBZesA1Tu4LToyaLYpn
3jh5gHuCM5AxSZ186dibedsES+EfXRYudLJwWU+TDFxXH1bC3jj41S5/LWMc/B3RnJPyzgZh/YWQ
EBNiQ0f89DPflOcPPM13+N8z1nSAC6UDwY1IXdmHHCQ7IMRq9CQweAWSFCBwfHfuq4oAc6y1hcyF
aUHk0vOusM6hU3oQ++E76jFdX3ZdqlQuoNSAUXQ9nSlXwABD9tWrNKCRy2GjCg+d+brmgYIM1TYp
ExaMUJV/pxWBQyr85Z/V/BtIIQGh8NU1hhd0UUojCJPyGBRFUxR2dikNPwbNH9EUZ9vPkqPsi130
dIo9c3i8L3qNl6uUPCglBM/4YZrvG8LhgUxVGoM0cPTOeHVJ6a7ZxQE1/MBtMSymeoWGQ6WXTWHs
/Gx6K4Wwln/boy9aeDo0ZYC8SCy6VU44pCWlaHMHAtzgGC3THn+FWASNTJJdu23zqeEGTKLhrOQ2
m6WxreoyYkiuoFksYRZpZVqdA40WJdtIC8vcKhdkOZ01R7/N88Nx7mstFKeV3eOof1qmJx/hDmSb
cTVndjiVbLyUmdLVGeTQK5xnqxevWk/M0UNAV8oNG60HeFYLSmVVIzrumAt1gLPQ3+n1zihPupqA
yL5jAI3Z9qrFvQPlrzTYBJKv4eXC83HXXl0+MozBw1rZTUVensKceutRmOE+7s5W8SP8E/YBp/aS
HWkEdrcneYkcmdRMeQzhjAbOIpzBCqASso6OA90fCVIdXDhhBEXTHuUQpu8B3XrRylzf/Mj1aWZ1
DmfTvGeQLq/IRqYL6JsspymTUhMreBRRIKxB1Z+CP+begCTxlkzvQwQ8kE0C8xGHs2KfGvmnYBMu
gcICBKv7gJ581FnCqSTT+s7C/U/Ib/Ee6P8i+MI7X7/+Vuyxu0AZ8qqUV2UglXukdokTFNf9O60J
Ys1u87oUFDOmTEnqjNbUHtqVJTSfDRhnEHkWAdwS91Dfp5Foy9D5yH9y2T5V3t0cgxL2C/+LXyum
XrepZr0DE7xKIKmOYEWWy1SmSBhcy4Ca2VBINecH+Xu7Z0gtyPBw+rxgswst7fojEKZyhCQ86gK3
o1Lu7WalTDKhKQas87qQeUodLY5H/SejQ6ZqC8/zEMO9fstYO6uds9S2seyN7rh53fkVmH+ikYYz
g4+oJHKyb+w/HVZ/Q+85qmxFPozkncZ+7aXHw6u3VjJlWezzzfgcEliP8LsHxYDOT9fcbPIAg0wx
n3EJ561GYsyLsrzCWl3L1FYTk17cEV0n+G4vqNq2iPatVI6KZE4XH0a00SC11hajrpOpd5pylwVm
A3aN7c2cUXF1PnVfBMbfTLwfsOCL8Wy21CovqN4j9rkcshfQIOVBcWhekMLQ14wV5uIUYtnLlBf/
R/DozWP72SPk7Mz2HpljScvi0dB9sJIwlXX/SX39A2r0yDSHrRqiKnSrJxEjt8KWR1RIQe919N1q
sLF1MdBcbP++IeCFcWUTHpo9nkeKjkktNSnpu6pbs9fQQcFlgxTlw4WaiahAav5LAorQZOpiMNYE
l9yF+ReYPzJUZ/+hzdINIjyIh5aUL1TJfGFj5nNsASptxWQbIdq9V5Loj8f2aS6WA2pK7VHdbDjT
F5T6oWKAEtpKaHnApFopaDXcLXcq28Z8E6Y3ouDGv8/oiwb9ZME1j3H8DZWF7Wpr2TpcRylqTIQI
fsoTCN0nskAn3IpfiaSmRrzA3+TqSXMSQd/Zm2yrfh0oosUVpzfnaflKM497hurdVgANMY9cWswY
7SOgA+tCEtt7Htk2+Wz3VYZolFLD+8lEL7vesrfufCbslPJksTHHMxBY6G++lv9l7UeJgARKGiwh
Ep6ToUWRt3RpeVL4Y3C9W4WXM/ixWx7vqlDPC6YLnP28QqSia0cIo4ETwHQJB84oIFfEH8BirwkP
y5CQoc060TXIysOmVX7fCrxla4N7SJlw7v3T6QAJUS+Hu1AgfBb63o2yGagLWI7JyThMJ5fD4llC
sXOqYMSrUddkLTJ6lf8/lx2+EG7Xg+4iGkVmm3R+dp1iMr+hRstUCfdwwiWgu3aBdTcRO15SoELQ
xHeUbVx1LkXFl+XbTs5FzxMu2wQ9EgZiRbc0Ik/b+wm8EglX81JEDupeOyIvKYmNCRqViaPaFact
b4gpC2gWdQDj083SG8EzjZen7+949kp4841Vi7p0B6Te4nBnQLCt+0cS5zYW806VhOPtJxTT79Yu
dJ5NdIgJgnbVmiLzkb6phvUMvLKLqNNe2X2wy0mgHw3HTvD1/4aeOg6SPnUMM85AkM8aC3epv7AD
bk194t/9CHf3cdxpOKuUi6uVJB4Evo4ah2l+AL4E0+/ElSFP/5JP410PJ9lSn9rBGurOSHYn9afw
ALWGkeLsFNv3lrWw0eaZ7K/awWVk4wXk9AvDrz9AP2y2eKa1NkwWb5bI7XHSScYIup14GoGvapGI
IB6FudKRVqPgS0GlCSeeqr3qEKsKw18wSwzME5O86tEpxujipPaMkZ/IQbLzGH+d5CeKnPMSb7tX
FZfE70lF1PfSQxb2vmp0inYTfvZfdZEUk2auwxRzBw662x+Zb/mt2v1AkpG0WrZuUUK0lSWtnzyJ
wryEF8RBH1tuxOgU5x7gusuzXDi+rJufqjdG4Qx9hKoTEu/0wX9zVCSh2Q9z14op6RsNFpyNdVzu
L7xw37aQyzCmcBgkkfGQ4e5yIpPdJTWgRdc8k99YawHFi2nPIgASn780ZLiTTxYVOHsTLJTdm4rZ
HO0pp9NOnJMTPFYV2HqKlIUNji4qIvFK2c/GgkgArdX80WPP9mXNaQ9I9qhU+byZ7dN9quF4aqY6
SNqG7ek+L5w0m0V534er5WuL+6sH3UP2MDsyAOjiNT7MaL8BqtJCeH1ACTdEzjffgf/ftYKLt/Od
Wnetjd4NtWWErdkkbdEYg5msvBzTv0eFz5rsmlTZUZMZtXmIj2uEMCtoIdhuTHmTXJPIGCm8tyaI
VGdL53lI719/ZL3cbQuAHV33QkJsW27TFeJx3jirCVYV9hLCONwPxnLdRVjd8Ea7hHLbXQi2m5jg
OP0yAZzFPpGvtmsZtVy4Qw35r9Ns75BeZhii8bwXjt+BcyXVWMlHbu32rXwm4m/fyioE3heQyuun
1bLicEZq0ZidLsA32LubfyN4iZNcSC6J2TxYwGV5ZUR1/mc0GF7As+jZS8Wm9dw9cu/t87aS33ud
gW6vlf1lvFNTsQU6Zk7TtaZSGt54m+/lDoE/hX7d7FQUnqWm3LSmwayTeds7mKFeKfiinqCZt+je
HbceiwOF/DFGJfkOvoNafDYAueCWBuFQ5+8hXR/3u57u6k8L/dp2HzBJaN5yNuI6KTggQ+a0t1cE
iWNP/Q3WeMEPtd9CI2DU23vDWjV/070p9LvWLVQeNXacqjmenQ8fleH1mPK4EpCv2LTsA0TMcMXB
LIBBAYgwD4vsutISF8l3luhmaEpRcJICNztNdFq7FU6ABKCdUZ8b+9IT9M38NZqDFcmu4cFHvVNt
PZm8lVVptP4z4n+3gl9geB+ssI8Gv5WwTKJ5M8F+0LYR7AUdHU+4wlBgIu6ICYssFynoizWCZi4+
rLCSVDXLfAxoPqP+9RElKC9c959gIFy84iFeungyMYlo7HFaHpFdvgFxwqaJkHENISHvrzOZUTBo
0dG5tRM7AcJltPTUId8TiiSmJvClP3nSBKgTfw2hVJINnfhZmqdIR3/MisRh/iwsCw3lFiHmoLcj
qlJ9CEn6eiBGh5+etUwGqh7lwXJb1vPUSwUpO16jsk4aQ0p1akIqsjp0C6RaxuAMWvGeANO4VZPc
p+W/DMxSFMt4iwKVX79WfUN+CT11wQfNtM3wS5BM4aHaSNPUKnUdjpW+q0oAtsZ/K2FKgVdHujB7
W6RwfTzYy2GYLqWkEI9+6GhfGAsZ17/1gyYIpDBu6HKaMcpOEToCb7yA9cAMljvzw/54Eg9FNFjN
xKGf4dQ1zoZ4E8mbeXQkF5m688n6EpNXCQaI1ZqbYDcTwj17la/TpNcMaHXWDbcnZm2/osU9H1rG
umUmKAnwIclvTZgrCfHRKTgVvvpss6R9fvf3TV9zT1fsgYPmjuY0rcBIEyBpCdZoHMN6a8BS6oef
yQK+R1GfL7Lg9tsyDzKqegABgaMtqJ5RNr1h5x58kkTN+ZPA66Qy2/HxsUGn94XLD+3M7F2U5uJO
/DxOyNVWjLWfQ4BDA8lhikJks4Yt6+j2coLoX8lDAzGolB8ClnqxbxdGWqFlZvRfXCKrtytZsY2+
wtAr7rJXS5JOGgSId6zAtgbHuLxkd8eXt3QNDsQ7f6c1QFsteUd0x45B3a9iHpPc+Xq5j7iu8HYO
0g9vJWtRT4augcDmINIYj88DEZD9S9bM4C2KGJYQ3CcIkyLx3lT1rkZs7RZ76xRUga7TH34tbbor
RQoS5T/AfMpPwyhH5SNVahWDJmwVvP0KoQ67Tzl0BMrXW9tJefWC6ohIduysxxNSW+snGNRWJrsf
S1aXEHDC+VUQi/RRNaqWX88cEbjRsoDgubaYQSx1uSkWu5rcGxvJFd9I9AibIuT81SgZznhhTyRP
yRwjB/u/l4+tnwwQzoeDdwW4iBoBr0aOaNsCkrUOKg6mswSIKyi3/TPCAUob9BojpL649fNIASae
DRPnbz1qc2pwkpd0D0qAdJjW022Z4d47N6rFa6hgcJmJEUwv2G9p6XACXcXzvzXSWpurKDRLxvL7
nEHXF+C2aZUJbNPRVEWOJXDgjrnGG/4WbyKxp9SMe5QH1a/t8S+kzJZrgyizzHJzd9ty/L5+nXpV
aROT2MkJqrcp0bW+ith2pPjWLdE8b5xIFOCMtGm5XygdOf+PThOfzM2vQ2/mXmi7oNzm5NJLcAsT
DRH8sgHZJaDwCCDNPH9BeqR5mUPvu/L4B77xhhEnn97+eueevpWh87Gj4M90Pbrbg07vqO9Bk7Pl
RpZkbbk3jYsxi6JTSOW/94/5Mmev3KRDV7lXK9j8lJVi2GSR4UjPNqcFJL8YbMMfx0qx43Mt3QV1
IPs3puwbSUcJ2cXmoAK0/E9vKZoFhAoz3ygMn9pJNA5YmPIm8JTMRba6uZnUWKMTnDRzuPDOTil3
FjQ44l76JumaQKiy1sBRXmbZBBejlNIFKNebg0kWIWWqYgEnS0DwUCnoeymGnsbbtTy2ndad9wyv
Iq8yl6ySCBssLpJ3vy5dO1irlq2VQEeZKUhAL9MB2nlrjFaZGgiEqvV2sIloJgb+mHLV6E5vz9GI
vI0YaTt8gVPYAtFhVQ1WhIY2vArt2TMFBTqI3OqIRYBnKtjjBbeEGPmU7zh/1ESskwtIL2B1TCNJ
21FDRBA/fHwUOrGnR0MWzsSbkeAfm5tL0SRmyhf9Y4qY1OjR8omAI76MgqbJqQG90diOdCsgzm/l
EbvEtyydwSoJAYyGOX/VfodgeItxSnltk3E3rX6/8wdXTmX+4uFxOpGEgooIE5/Xos+YjiE2Q8jp
Jk53VUX2qlIX+YwNZu0EekEvQGBndifGdTOndHMqSLQZyiVcSUTUbGyLzkO3VLziEU2u1adnXXKv
nBUKZh7MDmQ+M7loCt9Uiuu9brFB2svQ2SAh7n/sn1sfJ9JozG2od11FxOrzaV0eQlU/nJaBrkJo
ub+Tzu1yR/XCxpOhXSJ+W6bx4deor6ejYLJ7hGqCAGdtc1U10Spwwy+xNdM9QWOigcJe0sKtScFY
3TE7q5Qwjb29G4j37sbbBWOIU+Sjr2PxGmW8rdRGBBV7FC8CwO9qiszHzZVT4H8UmUdd6rmhOZcd
tyu9U9F02VN3uB2k9cChKC+7zQ6lY57TtDTnJcYmDjJrfbc+LTrudP1XxrsE0dDPIVSWDYAyn3sW
SzY40jXRAhOf8MfFz8ex6xtBKXk44zN2h94oOc5VItRYarUZq6ZDtd92t0Fh+9dNSmb46p+mQ+Qc
LsWfJHDSzSANLcAjXifMEgmbodoZNDcLFK56B12DiJYE8CCbcIXGCGuPq6Q8KR58icLcH7dVCQaJ
fdt3OtTkElBz/Q1qKV7H6t7/w4+6LoowrQzroGvUN1nik/Gc+u3y7laSVDutcTBlv4kBF0dJ5QLk
71ODCj0jU3VCkYJ0kXF2XR0zRYguQPsowYmv8ct79ANKIyoxhQt4UQBDD7pb2iEw3wp+H/5SxQYk
BmKTCeDL4mnU3uK/z/I9WqqH6M9ACw2Acd6PtJQHnAmF/uGrOUMChjFEK1kVrGwg743VUC7Lqb8l
vpe7Tj5gf9o1jxk0776LhF/VLtN9OkfvUac603yCYglyZyqxWPjNuaJH3JPqxzX+pSB6MTfs+sgo
SmAiYwS6qm+WnxMX/SFGVIDdjlN6p6QyzbGtOctxl8oBXyONHr44ulHBHSVWfjrHdHuI39F6swM2
ELNwd7emSrGXybdfDwiD3gbJb1kC0uWyh7jDo1MQKTKyS1dIMOPYNSiBLQf9f9RGIX3Midev2yhy
0OWaVluuchjh4WzTTzMV0ZJXzIbBZTFGWbsY2QmGbFwc0zaYvcZVhWWoSEV2aWlG/GiNHXPVZXl6
yAud/rSpvIC9I8zE8CJcYg8ZB1IwXMx6VS7I4IDebcmHmqZIxgj0mqqQEE7kxb4soY5/x/ao7i9N
Wq2UlZXDmA7GGuWwF8RAs/zzN1l046hVBIO7vcIxTlDjw2felgiXuxxOEMVAKZt+UdvNy8F0/6Ru
xyJAOG3munju6K1SIenwnqRLja7Ld+pfscRhOE7j7ZCkF3UfDPMm9NIqpKhu56+ZMw3hl0oEMg4U
Elp0O8416bzlbJ2ueqkasRyQM/7ORhj3osv5vI+Qxk1FNR590n/ipO1Qi1QGc82JpyfBU/9P5EDb
UDNEuX70fPk3OjosPnZuAGFm1/94vnqGQwSJWLcYlBi/aRFEmkDwVXq94Rg5VIrboopxJNh4X04M
e1DfMGwYecM3d4POK2oPDgY61fKbzHBupHOfuK6mnfY97NMjO6p9N8PgKVkq0mF23l2x13TEj5YB
OK0O1Qz4LWwGrQV2rWDm1tmGoYREeXuAHQ2dCyWGrU0rzqjjO3mQuldj7GCZRHUUHjtIEPK0oYhB
8TKatr9Bx4JOG7pn52QPhgJcFbCXsxBmcVbAUrcCA6vGIoIncE3bGcAlxD3ceKz9g/iKKVDEhsXM
cg9/gaFky1MmUZEFWbdrZbC6wVDhbSb5B2H8hA7KrOyWGTJA9t94rYYehbkjJ102z49wcYVCRPbM
M/vOxKB4+9vDzOUDkf9qU+57HCBQ9DFvujOz+1vIMAr/hah9L2IrElp16G5rcEh/xMs8Spaqnhsb
hQ3YtmcSU2jjcwhxssxR9eg6LafpL91Lk3OrVYeAHoa+KDck8rtxKWhqdbyDo4a+PeDadj2I9hdu
JhRRx0+pEWLiJrBYAIHQ9xWaxw9pWJbj4SwZFjd3QjUZeL7VHYW9QDuX+s1NyP0kkQx+O3LcKOvT
z5X7VPBE/tfZRhA9q6o5c4FhE2RZ+c2vP8AUNw64+pfjTDVykFJ8VjgFazfPtp3cGJmoMCMnZuf1
3Dv8mCgm87BnDVQtx48LaRgi6lZ+gvUrHOcApMl41wEaf1iDopBwpDV4KBBzcXxxSN67o9pDwDwc
i509Nu9D0dwn/p+mD62lNwbIYQAZxIjBz+Iw7mQPMA8eGJS8UmzgCY6n/pSNs5/b+l6TnplE0jpE
vMpszxmo4a37ZNd8fI0r3d0RgjVjV5Z9Jx8jm1YQ+h2pBso5JLvnLnY+MY/gAzom3ZPU2ZkoW7gM
cuOF5UzEPEuQQuJxTUGO/6bhjYtJmTZiIe6D+g/r8+wDvxb8qNlNW7vOjGYZJ/RtQNaQOn0WtGHt
GiOALn3pEl9HwgFNEBSPyvXJ2x3thw6ah5YNwyPgBZDcQdRrjyNiO8GquoXVXABnAVTGvOZb1/Xy
Vl791YUEE7eqAory+ixkEf4CF4rJV1kF7OxHUOAvCqYLhWxFR28hA7yP+RWS/4KY1tCsVzZIjkru
A2NwAM99wRIp6oTHPUFu92WKhlQNtykY3/VMy1H3WZWqzTgNyWHG2Pw0in1QkjRugMMhnjpgRUzW
GqUJQZifEimvo8HrqRfOw1CgOyh2+444Z1Sz7OelMORbfKIKsSGMsMNkhHjXK2SdebxK5CGwqY7k
QUQC17mfQUu0VMvn8RjiQyX5asROklmrcgOfCUWO8GirVAiuLernuyJz17Z/61F4HZfLhAq8eg9j
TaqQ4eBrskeCfb9LcKRd1S7c8Zrkp8wmJPw941WHIOSxn9zHaeNE9hfQziT5Wv1PTXcW97Le2LWx
yd8iGzCwXK++kxhQ9JUM/ilF16zQYLLIiJT6WRnFXVPs1dzQykKDK61MGD+Ew76RSPFG7afD2IZs
XqpHfvfxdU2EY9j78SPKyc4nlOab5ZQKs+8FxJK/GEuG4YRvP6kq107916Fxi5sqwvS07ASCu1bS
+ev1cTxZU7BKi9cxmF3zF01ExRweQQa7Et4PKzCusCKGtpXnznXDHzKisNSHIxL1qjUDp1UlK4p7
fmJqOoHKbbxthi78f5Nl/likIbFywkcObFOlxHMpOwJiNHbligJ1cB2Xb1PRcPOptvVJkkl1Xo4C
JbGxXGn3M1FDypERF/iE88ehkT5SY8Nhd1WtQj7lEOK8g9hFETZ2im08GfFIBLamVprioYHVnHZ1
WQZ9GkaT/toHHK6f7ZCoba7SDa0kGcYKTakEdOyRvvPJgIu0sWc9QS9sM49K+kYIZFgDryMmFVur
PnUCwW3K5Yn7/IUjW9jf98EjmA2eJGgWPIKy1AVy13UxYM198h56I+9TAgLKCXwPSOB4v0peUk6S
JUdLAarkcNadfrnZvun7wEXErVoYwk0lAUcd2ldnK8gI9p8lVSQTU3+m3o+I4UKfgux+1PcG6NrR
O4+38jx1EpZyWoWsEueupFqeLi7EYSWWeNIrM1lcDTFLcMSJPyzkJoEeeB1LIOjSekBD6yMVcMuT
z4CISA55DspmtwLXXgYP83NLbDcaT1BZawoa69nEnLxsHlW+zTaI8lJ2+YNmiSNBNYUtrFC5uGH/
G9YmatWCSPiNKtqhrHuPREJZhSPdb6bA5zY2dAWc5Uz+GPsdTm3dTXpaiy9jMmuC07L1xCFel0YX
x28/ZOB2+8YwaNrqnIfUBBr6oZcmscPJ6hiTe0fYuiW5BrOJDBj7O6JGjlyuWzt56cEc6LkQPcue
egeEP4p/jskc3WcncjVU+z73DS87OE11Vks+v5fHK/Y0eoqsPIkDzd/TunTskiYQ1e5i0no/WGsK
8828MUbWRiLkHKNC02n2fUTeRmX0XZSwVzyD/sVtYqDlaj3NsNLxzfmk1CiB2RHMmU0PyIZNK8p5
PajS/67YK/oKc7oebo+tjoCdu2Vz15+YSGsS3EUwBzE3MM0FGedOLT/NEkLDTqMC+Vo2ZNnJEB05
LXm7SZlsqJ6vsYQFRNq8PYxuTniJvGpHzJXDng5brXNRvQ0dwwcr/zhFOP+VL21e55Q1cmnwgIiJ
pzSTE4yhQWZyMq9tv2bgS+lEXjyQ73dbfOxSMFsNltDAbi2jo8MtFPNDsH/xpBCyp93qGavDY9L/
PgqYxUVlrzRON6+Or5gHyc9scB3XSAzwNCRJeQO4ViVwipkT2zvTF1dxaCO8mIXMjZlnbTMUFrJ6
fGBYNHQbTFuK1bxxT+enUEV7GErFfkNG6Q3Aqog+ycFJn1pepO0WEXziStduikpyXwHMLJLgrbAQ
K8UkpDTPRUaG2L94I6AkAln2ITCo4OkeA1aM+NLSnmMb8VaTtPxMgSl0WHXqN21tRByhxJKTLqtk
pBXcBK7OM8qfnNcnreGzPOupVQcc/WYiaycnvcZH65aEdLojqYVGbDI+IKBBMX3TB0lSofpoKPA3
PS8WLxhdGwN6d3peKpCpk2prdmtqrihFqp0pY237gvBHGdIaS9P1SeLRofHzLNxFFOyYjXFzTiY8
mj69h+1ESjkyKvaZZhr0Ls8qu/M4k8eFPWTsT0r/3QzbNs6lD4CDgQylO2NPc1RGsmieFLZ92/EG
ibUi3xpC8l4CKRNlYs4gN3gr+ZzKTzMfP984v6n9RQvzeaqMJuC/CiM5Xb1k6EUtU3ge1bIX9Xcx
LN2eDi4oEY2375jpt6kshw5ZCKtSl0qb6uLX1xM11uz5g+JXNlewC0GH5pks0G4L3bDb4RP/2cN6
qr8oVfjGIl4/xgFu5k/kPDgj2pXCqa0EgdJFMdb1P3aMX3SOsU8xqvU+DHSDycVDQbbHGmWXva6/
ii+yp3yb6ElRM9oTn0YUmXF2sX3ktmOc1Qm7AQnG4ToQyZr/iwu1yMlNVv1Kf9MIgPfKrIZghZ+K
RhloBOloxja6liTmWSWFV8RVev+Bjt6FSSV1n2GOZXrkqQyP4vDwfs6P6liCRPxGDXhMLxAuIVf5
GzW1U3k1ai08QYBAGls3b/sgcQJHD3AcbMoK3c4BLbCnKLKOYR0Kjm2WSy6j1pvOGTDgiwAPwYGv
TtYDUKFu9BrjIyX4AmJVW4Mfs8Z8QS0GjB51ZWl6pPZbheis/YWAP7RgvNYrZRXS/2nl5BSrreF3
YVLPolND7hrIsOyHFjZMzdalqb+dts1w0k5YEy8ER/ByGskq+kiFhMZYR98bixDAtf9KOHSlaLFp
tnC4/VcJEv6+aIq5VidPC8LOpqE1eHB8fKymMNqiyTFp2JDjFS6DuPC5joTlxdTIOLClRgBhwavl
e3zgMMaBXR5eQcsN929trtrb4P1JGya94pFX0pwi5jxRjjMhwqVH3W0XaDiyzVpt7Qj7mA7/nvql
ZSDXj4NZNJXJqlcC0XxnvxrBVPfmNC9FL3ZrEnEuHICh1JVH5QSTLZYZ3QBrPX2+94UFYI54vH2o
0TAd3gM/SGAsdMpRCaEFfv0oEVF9bMsBq3RqYeMempjWravb6UPiYt4sjyWQRVf7kRqds0iA+mIq
0XHEd4SH3Tvzfu8uNbkyHZA5g0g0QBFvysLpzRtP/6TxF5XC+BDM+n6VBvLdFTLdI5ykKjjONuM3
F6rcAlcXlmG69NydtGyxAvEvxKPLt4c/VZce+RMIgPVwdJTHmnFx+CgNRmdGa1CSafqCTyGbFkAp
iMp16/2SW75GArJ6F0YgF0LbHh+Q49bqJE0yLh1t+gIII/7sJCG7RwlWKXVDKbjPrfRl4pkVWYUg
KzjLFzlrQDbsGWZxUucmhpoSKHErFcHag24KlBCOhihzuQyvrbZ78uO5I9YC0q9c00VFrWdIO48U
TvM2X7hk3Ja2InOQ9jvG+NrRf6cB+9D4nwPy/wz4rnH8o5YlPwr08bZKrai3/cuQbbWvUERG8HGK
DytKX9rKrmG8lQrfg8tN8REelKyH83gaDCjBm4K45V/v10aKd2zjS6ZKvlmap8kK/lB8ZzkuVHqK
BzPD/TX67+eyYluUyBiMndpks5Dr8dgCq82NQwmI5+2oBzZM1bWQoVklhKjeUpGmZaghR/tGJkC8
m4lqaxA9pIndz1In295607VU4iG8tzek+VfLQ7W5VHEf9MllngDT4o5LITU9k20qlo3inhv0G/+X
VHGlwEGbyM262AMDGVBDDFi4CsrVs1B6vqnsA7e01F5b5anZw6xgL/8mlItU2Iy77XQLUmxaB6Ak
lYhKuZo6GKxs2MU7BttkqaQUaFWJF4xwdRdP1N3Ukbj0+ttUs5VmFwiC5pTK7VXlvfcEFNmnCnpU
5VlXcjKoRXEeoUMUxnZW3b92fT51FsYfXxY7J/i/cUILFyLR/XM2Slu1lTeYg09khfx29VBnY6A6
ZoKGoxG/SdkO3XH/MuY5yCoOfxpPycEF/jwCvslhlHoPPNbrM5uXs4gyev3IE1XnZCecDHWAC2b7
GA7ojg01hTvSlUQCqm57bIEzjBHgFLhL11rsWHqSP4BHakvKNJgCQd7jcvChDkOanm5I28PSpZAJ
cE/0SfJpFrI2XhnLfzVM/a9aLoLCddrbFcho3fp6NPSSoWHIalCyoOOixeOy+G82xKqpnK2hWLKm
Jw05n+utZ6uDWeV/jkJLl70NzEjF4sZgGCbfqH/OE3MjwfJ4nbXYq7zTeNAWL7h7o2ADPdedA8bw
n8p054USjaZRbz9h2uUf4OIiXjEshlToYMLm07oSqpcFntLlbFggqH5SlR8E3jKGpBASJHIJpQV0
V5/N2LQh9SpZKW6cBijHVG8qsxZmIJU5sVbvGdjMI3KiX1Jktt1ljoXb+m4odRAO08n5nk7rb8ZD
pa18wxSIxXApSnn6KRKs69WNUq4CrTpUqmf7hyIZPtF90RauTJYQZoA874BmoTltZp1Q6ENZI39s
8mkoKZr9QQsvtR0Bsu8zI19pAAY3/iuvo94a4yrSKxUTLTeNZfAwtDN9JfSVzXeMYCCApZH5Vpeg
lXQGrdC4rdezmKzmB5k7cDdtrrDZht7rCxWnsEEnpmrXrVCHfrIcpdDI/6TfpbZDdewl28YGltYo
OiaIozN4Tg4uGJD8q5OmcnEbDyuxrHtoGViSDaLrBqRv1Bz2O43IfmyI22EdX3BBzyTBukZA+R8V
C4USSSLJ+xTsL8eJwDbJcCkBLkxYnHiF0aHzGJ090SgA3e7xxUEslQYpcKOd3ksxEdOeYxAjfmfp
wTkfg5T0GhcJFlKyL96nA7+yKPVMN65fgk4AUUqdU4CZrUVAQoRK/iBmMYm37cEyFH0V8BHBljx2
z4mdCSgJ4yAa8P8TWvEjnjGss9hHnW0dVxdeYUnXdVo4twUyflz3AkAKwU6TTcF1c/Z2RYGJuK4U
mti05OD2HOA3sGmsNSNKqSbNLHM6JJIxDoC5W8H/EAtUdgjkR4IXk9b/PteVv/d6W7P1umyElzhv
x2k4y/iKDd9DJhBRxo3U9cQVO39tLN8KrJZt8MKG3NjcbFWto4aUBhwtXgO/mj2nva2IjqCip9wC
fQOAIKBzbwn+1low0IkWyrgvOTB7EN345yBnxteS6ETf7+0Adgovc058ENiOMFZbAizJvruokjVd
vixeCA+3w1D4lfgt8FvqCOHAHVDeEMrqRBVaugtQ2N1nWwL5NyJWXsNGEstGQiCb5M+M7w8x4JGb
gkm9CZm44iNXVbpOadWUqzwTJi21lKA0wc7BluPMDU52rOwVkfYGxqZuv3gV+tPSnEnRPzPpXQDu
qXytonLptWip7g4EoA/CLzid3Tos84Kdk3bMCLZDT5zp+T8Q0p4kO+aLhx3M9uyP/NqqVVttjYyY
QhSNmcj0fXEFpUhLAlrdc6UsAWCimBUgcBRhhlRgoaKhpdPz8j718tvn3oXRWtOm9jM3E4MiyfIp
hipnRa09DO/KGnSaiHENOp6hCIe1Ge+3LVKsiWBGfT2WuRYQ8PgCbuekl6zct6NR5bF8Quu+HjKg
WlWrGAzRTnOYPBV0d0Kq95rCNs9nq72gbTUA4ZoE6WjyDsOUw7SzUdPe4KAWFqgyNfQg7bMCK5AV
UdveY7v9IyN/xpNanvlIsq5JDI4O45VA/WQOn4uEmZXLcMkGBxcjstiMprmK0KS5AKCNlzY/yk9q
WoLiPc7Hq4zE/BKiVpSz/7L588qmS1ShxpneRZ1AZLDhSrzJgiQUXO8bqCwwn1tx29j4WsR8wUtb
Yc21SSpAE1GJYVJY20oQ/cAJqQTQWRv5QzkxLPBzBTpt6V878iF41ftjRGR7sQ/GQn950jZrrYeO
ioWHi4CFtaxaFN6knE6bMDEexej+Her0i40OIGf70pxuZgy2roSw7JEdgFmRvXfO3RE2aUuOYl4G
rgPk6JdCCUnoeZt0/eTUYbXYPM4mf3H8F8les/Zbq4bo+Gs2fXuTTWQfK767cGdfWTkb0fzodYCp
qB/g+idpOKETaAD3r9noBDitMXQUwcre3hD2vmFkzZVDDfnyhWxFLp/ffNZRNdqg9XKPAlbA4jfm
kP5JmB6WIq3fCcZoGtMoiXIo1s1BMPUEvgAYlMeXuzAOz/InfW4+ZFSl/AIK24jEwZ6Uiw9Czvs2
xzoAbZBZ6qvjUKP8UAxyJjMipRgcF39lpPYt0x9DyT/NLAuE3XLI3dpilnz4tYvQSpwbIwk6zrae
jYJqdOqytd54bEAQWt7hj3+nUkfeE0QzlLpDxeC4nMJR8ztRQ9spDEKOOSpxlKpBkdN3II+CyKDB
xQAcTUwK0ejcBcM7fgFzB5FiQd2/f7slT7rSnClmjexumwnFcMopRtfnH22maEWCHpAjdpeve3yq
e+Cc9G+5UvCfaxFQhqgKGByRaymC1jYeR9Sh4bFh2ZBVLgwbe/KerSo8TFK2UBUPnLjOcechME2f
XImuCniaQpVxq03C3rz/5/1YmT7HPN7E2X6112XBCyPY1mg414p4IFbpTHJPZMtN2PUe2Lh4Dzbs
FCb9cFTN8P4Qk95Q0yzCgUISxAQ3apQmHKP025M9cASCZPQa/+FQmnf6NCXsH7cukzgMlxLWzw/R
FD1s0uuRKpUAdHNQV9e7l6LisRcxczBCAjirTho0HdwpwrUb9C1wXmJlESkY2DZVVDH2pp93/BUO
mmIUySkPp00m1K9z+Wr9D6FPlsiPjoNafJ5pySSGectKDOu51O/94l+EKSVxoT9VEmYp70RdOW6N
2TMJck1vn2fIkkb+uOqPgmFYeHEWXJwgjbgIftnUSaAwEeK+4hnldMK5J4QK2v3lFUT9uhy9fpO3
0D62FUAsxaWeqsp6qahNlStyJwEieVAlVXnV9LcbLoN/hTOfPVoR7tWBYM2BtCwFu90Xo2cJCCfx
PXEOcNizgLCyZ9cMwnn/Ml73hGwWybuCTJarkKMNZYv/w1ql6d6Tjj9IwgFB1jTo88ME34407wdZ
RSunZcqpMTbMhuCt25AfOYQ0ixhxSW2JWTAXtRmUir3s5tKliZzke507FH2tVDa2pmYy6OlXme+L
VjnBxJo8U6p4hMPZzkasdV7grk+SI4c23CpEX3f/kxIWxiz1p2y8vZAVvqI6ijJCseR2eyNldaCH
jHGy37JUMmcjWZl4Y8RavMC1k+qYdUhpKiWNiALIy86ffgX9dCnB85Z3gX8MvL5TJrb6jpJi3sEj
1bD/sU0OCHRU/jBcQzDKWIWEIFMW+7MdyPLxTcGew9ypoyR/QIlQJeYPPFXO9z5c0UEbun1+OeZp
4xVwm0Ke8AHF6dZHu/1bEjL2pxmv0t8hLLbZGAof2yk/B2E3/QIhhNEfHW7347GESo93W4x73pgN
rYrE2eRhxozKYulLIG81HNqh8jWrTIiF+/LiLAp6itpePKPf2OU23y93NhUsMG7TgpFTvg6J5W9m
xs6xVcbx8d09DWLd+3bYO4hnceg/6Ghi7rdNsg5PphSjweHeQYoOKGPAv2Mqo2gL6Nx8lx6rjYvZ
K1Fmo0moIUQDL8EM1h/IPdUIVdb+n2SqeR5SKjhT0H71Y1qejjPjAeczIXJca97O/nV0YLrkyFoQ
cfsKevy5lh2BLSHqVzrWNmQ65EdGMU1ki7US6rk4O4bWBpv+gNM9HdoQ/lz9AxtnNA/gMDcaZQZ1
PvEMgj9XUARvlKPfhS27sqogZORJjLyN7LQgRqm8fYA3AVfTdUnQhvZylpuXyC5/0JZoyrAddlLV
GMZttBzXP4Xsn0x3ut3hS4f3zgOEJ4h+ARIJbIr/eFhgYfWh6oGmU10NsUTMiOyncPkdPuyTdp5q
6kSsxhtLj6rBG2x7/TVEZ/5tDliWFQwLp1hjSe5+Nl+n/5wZtmB7JsY9LdRj4ndQSTZ67JWSLgZ6
dV3xMOg8zsRQC+PDg6/YX7NE6jfadQ/BI0/fiFN1QvbE49+7WWfrdXrSIMYTCGxF3Cta0oKEh4Cd
Cfg8ZVb+NQ6mmlD3LwMADBK47XE3bS/v5gS0MA/w/vBjhWhOO1tDF0/LqMs5DkOyBivdN+lcPuYx
wgcY/d3Cg/fgo7CJxNLp/FliZf2GFuRDMl+F2HlCaPf/7fpX8XLTBi0OPffc8fFMyokyXz4V8Gef
9hvI8AmlaU0H4sQeEejlEQOmtjD4gC9lPg38STxH4Bkoj4sRescZMk/d/hMeysAXDVN3Kpx0LKwv
afqTbPksAEpIHbyQisxv+c1u6UYE5TCamRvmjw7BZIixza0Rd33Nq8wZpOsOqyrEvGx+FLwYsLkJ
5QtIND1RIV9/A17hjzjgdbSKB5Db2kHAdtttvkwj1uGLrPnA/Gn3x3ssk3BMhMv8Lv4vohdABOcT
xryfX7V8TlQh8mF0By44/Jv6xRHm8jq8DREX0GVbErHvUWPoeTmaiBCZNccLdiTE1lLdv1mCTR2t
8Cj+I4VxeJJk7khBgtlv6/Tt/3f1AB/eUfjxPkSTcVwyuStBD8SQbEJ53Ksrkpv73L8IEIBTKNgz
qxAiwZzXbwu5Vdf3vTh0rUUBkC7pH5Il1dSJnpvD6U8qqTFR8xJJV1dih8uu+HYvsf6KQcl0sc57
E9zBmGlimmdKu6JYzIqQySuPCxKerZs43ZXhRbPILYCYm0ESHncyU2dCDgZG88zBpIKjVlSuKAVi
gcKoeYiUL5Q/ggfRFHcEWp+JP9kQwNB6JYrqxAqsq7xNj73VbzX9abaRn4tn6BkafnO9eswCMO0D
psNiI3HURZM4Th/bt/RkGCeu7LY2doMVYvvdbrRvdodYcNv+O0UL+f+DvXuDpYT40FPvTIsSXhbB
DptHf6bdWzGZ38Wd+Qi5/GetW6MvYneOThpfYn1cvrxcJ2g/PDp8qMEEY6FBs54BXqYCo6+e8spD
Rq5br8hPpbaewrR2/OnM99rG4XVYVgzphqlprKnQGjNLogxrRNOBoVMaS1tENJAEBvHFEZzX26aI
m0PD2Ycfo5eDcBsNcF/hvkSg5NtC4Q/gDSmCu6rpFDlJdgaQiROCipgerbuDKEBvxJUBzKkfSDb3
LchXJ07EQb5Ax/DF/7JZGKumHKDGRZGGdKbBzy76RpKCwQoZ1cbPMS7ugzMiMg8Zu77EyTCYs27C
Z4O62n8aLRdW43WxLim7/QiqQ8zBuRXnGogxkjyVgGMeGH42k6diOiyGVX6w3DEjMIha+UmvM+ND
mUp2EoEOb08V4L5zdELFxejQerlG6c/91IuXlyidEYcCgf5C53bb0xBObeav7eptZWtfHfzid02T
lTDHBmP5GqAqMcsyzEKxV05Ri0LRDnLQzML4G7oJFazVEPl5o74X9ATP2BBATliDow5lSjK7lsgd
VCXq5Nk1ZzCE0NtqaMHZQVcW5v/ysWQXcKm+G3JErbU5cQGKaWN5/x8SiZRrEVkvpKmqC2jNpJMW
ZEANeGS8bdYzU7Z+6bZEaNrBSQaI2F6Zj3JXXQ//JuISI3aoQgIM6PEETg6mwmegahsSpa1Ilaoe
2fu46bcGZrbFbtLAVa5O/TXHgpM6TXW/dhMS1BNMlQXYEqNtULXjSrRcz161jWCvjzDqoxbwHu5a
gC0SVKu1X1CWIoFNik0x0aublD4ENBJClOCItXxPuFGX69JKaAYZNLLb+QT7IKNRxt+khRFKyHRr
ZjlG0bOsHvv4f+HXmr2W+rDh+WYR9P5w6DejHRbBDWM04BRV020n68caEGmf++eRXANeUYqra+pg
KlR2JVHIA0zCVgEDCjasR7rYwe5jvHuttb0yI7K0AN4xhEjkHQaQeZq7UkG+OoN/n6fP0Rw9fR8M
f1jk/Zezon2xtJAXt8oltSpn4HuSx9yYTkra4vwR3vqPvzuDNp6p1Mtk3G9ap392KhtyK/Ug6osv
dEjZcTOe/flW4VRwJJM0D+36WvUwISgVcfwCG6xOfSqe8wMj+RWJkSVOPpApmLlXVUb4vJrr6d57
Rl2EcfYH7n2mXLaLjRLSDxZBuuiaT3DNtvl+M05GUqgm/CHobXE7hC0rijTViM93ec3sdkH3x3MD
sTTjU50ARwvrMTeNiykfCTIdnxwv5Hvsvn14mPlN/GcDH+eJlw9h1sQKi3Ryl3/XJREz2yeAmRuH
5u0U0RF6bFdGbUFMqslE7hEWWTPbD1J4bkztyABHniB25X2XLrZ4YhfiVSzKyMyGnU6Tz+l1wiiE
SCmChrVEPhIbJRfzknCegZ3pwyqo1KCklnUOocqCDr1UkXK0DVR5JGILatZEwfZm4Z+xaRT2jt1y
9JRbzicInLc5bbjwzcrRgt3TCohk7OztrdjWx42cXJO6HbDx0OP8VskQw4uEQ4/DuirYBp/7FdPQ
7Kk2XSemR7wS5FePjLac8TZ9nr1ElffEBPoOP781Qlb5atwfa/CfURzchSWgLvHUXQ8JCem6+6zP
swBqbvz+fhqCVR+BNe9v61VBTuh+9OkG4BOlfE15k8aopSB19vDqcxWhxS09v/8S5ctEM65F09rE
hGJi/dNIKk7UQQenDq29qvuHQVKBA/I+xTrdxSTcEPE3oyqCKQBEqfJ1COytuaSoZlKgKpystgFe
cH7yZE+2oCyW0pr9dKNUKqwiUnXdGFBfQDOd1u17OaY/MJsdspZzDR7kSvj6VLvrMD/uDixUA+KK
7m6mPowONOWjII9bC0bfjHI9xWWEBlreLg6mb1UR0uruikpy6iWJ3gePOL4LcA2H+KPSon6WpJN2
0TdHh3y7YAFUBCA0aP/r8N0vWnNqvGDgllZcYiesdvxF/zNM4mXlT0DWEANd7qExSqeR3bO58k2p
XgIqmMWWxK7D3+Gz3mpnoM9AFVFvFVuDaeReLl4go8bE+UWKonLhmSfNf3K3rJIaPYlwi5dSO/3b
OWppqaZDj9YjIHR7jGs9aKeYkJ3TcaVy2Rx0DOuTX7hbuNIBnwOLmdB0JOQ7hprfcVWyriFV3jo+
JVESCBKJLHjr/M/e2BJhh9vmJcAMPT8aFsUlHikUK18QEs9kzDrGPI82vbd0/qHHuqe2Tp2jfmFr
C0kqL9lwH9rlXsGg7gpDXx/2DqU/+BUjraGjaDJoS6M8ms2CVuql4EedS4q9YKCIuMgwaKHIAAzN
S4oNktjanRtec7NuhLJqNrJp6HsiBFAdMSKFwrombDnhANubV0ZCZOcBp8SaM0OWFhRwvHcS3LOs
CPiqBE0WI11bIIMenQgpJXHL4VrEF4HnlGQP0ntUydflQS6l/CaEl0P013zs10G6sa+27Rh9bB7V
d3b9aNiYx/KS5EjQDGK1p2I+eGCsfDdvKATzWZ9TdDCE+ss+wRBIPfuy/q6PGLsdOBi3UloAFtHn
DQ2N6y8MGDwzFwZmi9pJ3L+L/luFq7l0tXr75uZz3xwURUs1joPRp65nsFVZkXmI8dHM1wSovw3l
hN+hzZ/bKXajP+fiXTvXplteB1ZBJviIOVluyQUgrcrDEP0xnVXzXbYWTKUB+iMRdq+y2lkH+d4Q
Ov/rVXVnbg7o3Y8wCWIwYk1AvQJLlKSLJEDaa8OESaRjolh6VW4N/XzmqmjhKkBHKtgNM6Leb2x8
G7D0oDEsMuBqKe3bfo0Ns/Rej6wz6ojnp3wNwzzy+L5nhh1XecDsfpYnrfbCYjM/NLQUH44g47WK
QsAMe7Dy3yznuMrktfiVijscaiVPqk8L4Bw8SU8tJGsw4Z1dj5F/Y6aev8IAFz1umUikbNGaelR5
C4qbV5cKquLcxRUrDahSVDqNX2g9vCr8nYKwvCtyC9Yx6GUed9KMTlEaTR9+gFXBXs1tTmkX5Fc1
lP/hnZ1fey1UT7nrKabh272KMEW6+S2asBY+URaz52/WlN/n5RsjvgTx1ZQqnrD06I6paN/esaT7
MCt7/HiffICnMOxtnGYzFbq4cnGr+qxsrla/jt4eahJOkPc4kqb6uDrWUSIDYHTs+B+t1+BdGGbS
8m8GctB7tdm4FDWm20npaNXvPiKq/wy4PFpVtoP0c/+7NbbQMiSaXyKPFn5OP5kcwxunSE34V+r1
vUBCKwabtW3yjyKSXrxCpWcfmD1MDfmBm0VMVUhY4B35jokCziXFNpSUIAg0uZPLD0dYbkanUWL7
PrZpgwTt4eRI8KCRTIs9b252Y8g+wDOc9V/eBo7tfz2vxdMZnFU+Z7uzyb+r/ugdpoblcpGubnJC
oZd68YmEgUfAtsSI3ZXoWC1Ujk2SsHAh489IvBfiTvLoECFfKdUpyHCrJNkp9AHI0v8JtGlveuQ/
T1fl6NrijRRVldNZhkrciHKwZaeqt9dLKf7PywLrtdqa5LAr3oYYU8vW03PQmPaHjjzUajsD6vMR
CSP0OsMcw3RCI2wdtnwcdLcCX0VF8XKjDFefh6puTQ3GUCJviq9AvZEM5z1MeE6V0QKe2EMGoq3i
xdpCCK1qfXMMy0tIPg5u8uBFNOQzQaaUAaNIznHeBhzj5UWf1YFGqpx0dJhOP0ox38DQYJkWkerb
nVatL+gQislab1X0HP2TSWX3ZnmbHoWHuZodstoaKPMd7R1PJP/snp/JfVJIvz8MXUQIHHNhXDZE
gHVKde6oKW/trWNi41ttyznuikcuyiu7szAXHP1fx4leT5Jvkaez0k2PDLksNj8PAgRAyfI3U1GX
dku5Dafz2dS5RwMlv/Ey4qiKnR3Lm7KtgneO5QHUrBfVkDq7MhVSrI+g7AxpcAJqwxd46S5kAQHr
weWICEP3MgMrgpR1ShsWkLO16ydSKOIXO0YWuc8P3+eDqrzxIRMDZe14zHwYKyPWu8lN+whsKabi
D7QUCIhpZrEqKKQT7CYusTLHHs2aoaiGGRdVJguD68IyVf2DrCRi9IEKUWMg7sP0lCyvVmne5NOg
eRj63rvkCS76e42nieXAh7PZAY6ttOc5jpqIzLme5yNkZKitdqeVMG9MrK8oqLPwnNg3okPv9ZDD
mDjKHvzJqCurcBY4IwgeVkZfuG1lcQN61vDxA20MCZklTMqm9dMt4vJL0XWgs0cTplEnRaSPA4Fg
uRYNpg0nmPYcsZ/WSwT6dU/eeu3y1cDv62yMl0WDxXh2QmzVlzN//n1P1rUhex/cEq3bWI5dvUnd
bxlTpSSF5/ErqY5nQeU92FXlpmKVjnbKB3xS80iceZpcn9ePJWM7ZQ12od1YByfvtBrCUNQp6eBf
TOi0hSC1pK3ZBQ8In5a77OCtYTrPBrlpx959u760m1kSW35gG/wG45vrlkC25oVIJEfv1c+GbiWL
NLJw0EYG4vcGbFiSOvygVKaDCKm02yfG9HGVvARtfyQvWQZogJpKV1BpLniA4u2Uo4ghnCC3+8xF
1XoSOOZSyHuMz1jmIRIVyHEM8R6ELf0dwDC6zuP7T66nGEmQFYagioCyYHPWbdOACkMBGoXFBUpo
0DNvDW8KNIjzDJFKChHQnysAo9JUxXLhF/2OntBrrf+3/WpJBJUoeJyJHzt8IhWk1GgME5YJ7AXv
z51rB8ThbFkwUC0N+L4FVhfUub1Bp5seXlcSStq1QG41S5OLbHu1vkbwY74knkwFc/SXVcP0PURA
rCDWa/r2Sg8HxJfbLkAkKohU60yX2F7FoGxygehVnRBCmjBpNH13YfZWpC3YDWXmYh3rapH7oxug
H2uKDR/hdqG4tgKQs85C64jZFIuaO5KINW5XNo5RiPDrctTsvzJhIdC3Uoc8OL/KJXqJXNbFlHF0
Vl7guiUrai4T0atYu61rubmo7te7iQMVQbSzuh70r6ap1CURkVJnRLylJDliuvAFmN+xXa51rI5D
Arpya1MCDFFUatvPXHFh+Ma+yCMfTRmTTWCuLbUiKDz6+ZPjxHW6a4gt9vOnaNmp+NXbP9QwZ+NK
DS0aX4pPuZJrbR5x9UVBVv15medY6EnSm9AcijuuaUEz+bkdw0dSF6M9qwQHXXRg8mxbOFUQqjzS
CAifsohFkCUorhg921sj72h8yMmC191F24g+6C9EctZaRIciLA2IPTP58NpVnf/VajaC5Awk7B9O
IZBVXhrUd7O3+V4vPRCCpfWM+P6XW4WYW8fNOo9z1sSZ2bDsg16mVy7868V4psyDFLExt8FJO1/M
qpn9jO3oxmkQl7t0kIS/oh+AuCH11GCHArOvIzqf2NtO+8qRD3i2+UiIvykCQcimIPMECwNQmIEC
nCwVSdJnUHD25c5bBrS6laoZSQMfUFaOX3jvnRjoYmwktHWQlMdm/FbUZ5RtNE0BF58sk4hEXi9G
lZeXgdMfy1LmCLOIYOtZh/Uz4A8h9YuMCNuYyU5l5Po+nG+0qj+qw9Efn3Yx+FRr33FtMWOrAll6
HQtBxh9ddknceO9JBHIyK5VsEVm8rMoMKQtsh30OFgXrYPEPHEHHutPsrfR5ieOsMvDv2BLLX0W7
3K+n4O6cAQMxum7vLprzJqeN5Np2sTCKJ0zA0UpJMZUCslWkFmvoC4UeQjfsGD+m5Ko8a0WctXgN
EmwBkXEpazF/C6OlQqSRf08KdffVEOWC0ekFvhs0OuY8RPHJ1u6N00Qt+vRt+7zOMHoQpWg/UuRO
oLQ+pU0/XXeprfbHG+Dv+GdgRRpjoceoRWX8IGiwNMuzkaEERETs9/zTdBYLgPjmIDsDJ+MGuMUL
bc7XuEJix9/AORDy88P42w7Cx38WwPePB97upKxruIZ1h6eMw/AdC+XEF0rImelf2Y1ZJ2pIgfIt
UBicG1NoIoY853yhtKnNXLi/qR4bY0/xWXb1H1GuZqqcmpNmXmUgkJ6LM1vLw3mteXf2esJRRNie
eyQVb+PvnYtXvtxbPkwlQhb35l7/dzFCDNB9jjStTtGk+xuiwIRajbPvo6Je6jCPIAcASSBcK+B3
1sqVURkk1sRz3rhhtSkAQWfOLN+0YzFeDXqkUKWAmWOsOtX9R0CBcEG/+KFHS+GMiogdUMgqVV2R
eSn4j1x8aDoNHDtL3H5zSFOAwkXxayhBDsbkF/0WHKg0N0xftrVcHnyYiPirERKn0xvemR8+F4YE
11g+AConPAHlxLAkrz1hbMD3JSDE2aUTN5AWKQvOjIYOo1kgPB+fFb0WKtmr/wmKFoOUEpeYe6yy
R08mc412TmKZMEDNBt9x3I+SOqMa1mTKj7Yeeujr+srNwOl6C/Yv8PiCN4aSv1yB4VXOUM1r5krF
OdI3uUiLk8IBHTuOAUGaKPBZFW1qeox2vht3mvGXM4V+jL8WIkX61+FQBuHoSFQIUttf04Yd8OLb
Vx3sPMIsAgLH34mjzcGw6OPvXZhpNzLM7yPQ5qxDcWptm8RdF472a+WtWz4eocdSANREXDpE5S74
rHVhsOkxiCd3lV3Hw1J4cN1hQKsJXY+vvpHDtRufwLUYAungRJcR+NvwuHhMKg/5+yD/zFp7Mj47
nmbxA3xTKO1LfP/hMVW7alkojBX7BzhT6KcM6v7u87rucspZXCya5kUjKfyHImx2WpwvfQ+ahtxd
j02lKwoacz5CVpYqzgFhhFCmtfZEmPX1hzqTxsbceH7DXGmog2nxajkELg4sZz41VeI2CD330Xag
BiRN7V7lZvVuc5eq0+WYhYeOB5dgPfHnQyACqzpQh8lSIV4fbj7/hZdRbURkC4+aICuKMi49SMCw
d1qXm4BStII6hj+RPtjW4RWtOzCnCL9wvgBXzFTSbhFSUXEbsaNSMCo5L0+32BtcUpV9Vcq+6FNt
qdVjgKwHzQAgAl4uekRdJjvhATpqP5VoRyTrb/cPQa8XpJC0MXXztyv1YlIcTyImjhCh78uFw59D
OTrSGNmMNAVEO/qcq6WmPIv9joTgoCWznO4NrFs7KFdof3Lq7kcA3lTNfu9N1+UdzRJhIXOVhOaA
QhRKDeqMybNpZJh1qB2BF5myU992lYMd3IGKdBGltO/j2xnuygrYU1kcoBMCNq9yIhN+AyjknBQc
r6Masj726q6vxheRi5n95wN8xae/Cha4BJ48eBbiTONrLF4IlIk3AI5vsHmzlUVjPBvO0Pcnm9ph
fum2QA1pdZmAgfvx4R9Yj2n4b7+UDoKXIOmhFYobnhuq+CUSJJRSpQmIXqpvabY8LtZtpU72VUih
buPcYHTEA9sV9ljRH4wCc/co1j8LBQSGxNw9RgTMkm9dQIjNF2k2MxyOAEcQWLt2WErpKCTSvK/m
VFG3Fpwl+fNC/+dCpG/RkaczrixBAukCaSrwSv4vM6o2V207Jf4o7e0K+rQQSAm/eXdU3m9wo6Dh
fhvys+A/ZqMKJE9YLg1SMpD3hzCKSQj52ORqpf2aoGZeeYeCG/kPHVED8E2YiJy5UobwzVk3dg1q
EHE6heQWzM2Hvn1bhwjaE380wys2R0p3BuqretFfd+xUMTMvX7a6q+8LwtT5BTuR+hBNTY//53BX
PUL5l9KfWYVL/iCVjVIgELwvLRxq3ZVttev9fi5XlAXql1YXKDndcsKXPdXqqJbV1jNzKXUpv1jL
hjtmi8XxcLZJ1HVbsLHAPO+L/H/PtVge80PJI5TS5Yh+bRJGGb8OEExhuyk9HHz8wU2WyhSwbrMz
GDKVuoj2v+O8n+ftutXamiUNoM4AjLDHoTFTm9hoCgr12CgQ2cZ2pwg54cbv7EWaCXjhPslKOclF
RYAfES1rq+sJuTcXtoA6HxGX9+4BYEXwo7mxqAk13XC7U31TPD2ok8i4d/73VlA269+Bf6yKb7Rf
+q9PhGDv0SsHPAEO41R4HN1kDXuPJPls7LquxQ8WKe1KoRtgPvFTY0KqugekfuJ6Cd8IXyLV2fa4
9Z1SyXmOjEM3DtpYj51K4afr67jT1EeXOS8WF1tjdN1zqmCWU7fbzn+zqktZKpb2l4Pi7/j49kb/
R3yd7Q98BbLRlsh10Q6eiCs/PHlppCStMf8bOR/6HWwJ2oLaYb4hE/ZcO+8jKbdJPyoYQHGpkocg
2TokESSrX/+ZJ+IkWYMTdv+PPsHt1A053dfBgv9qgSjUD6jRFo2p6pmOfGRhvMNQrgtbaHn6bhlA
H6yJ+PB8XMnY/g/WqnDRU9ZtwSUeWbZryLVtipWnwz8uzAj1BZgTkvwrrhOX9tDsq2ruiSgbghZb
CN82XCUZMmWVIUO2y5h4pFTkIPh/tW/W4QvyRDNFiPWdWPftcPBNYAR8T/AnAf9SYuvVE3Vu98zL
7WVOAzr/xdintQa+ZIUQ5XqHXNdTsXqr4gXdd16LBM9TDq/vBMid4bpCyP1hxvttuSiHFLu08zFq
R2TkPXSbgNXzJbUlH6soj1hQ+dzrmlCDmFciD/KZOwTqi4m2nFn6ciOvRUUxhlojLCWjwWhyndBd
KtV8MJWLuiZLzAODnXnWZatw8KokS5ymONDB5Lf4JSNIJqK8VLO7MJ3QX/B3QMWsCj4OFqz0KVNa
mjM9aM/GtwDWr97IA2OraPGlX6rrYSRVwatSU6d4LC7ueKEBJG5Hz54taax+AVLHHkOFMLwaAh/z
bpw4lWUpTOivkae/V+U7VT1JsVuPtygAPH28gcz9BHPT0H/5kkT4TXxgZ7uwZj/Rj756yYcRoygy
UPROkp4IVRr9QcT9iyKAepnr2rs0/+z6uzOj4298Z+GuUU+y3LSCrVVaS/BZy0uAXR8Sit8Dbe9+
dzj9S2MgEtLxgRglV25/O5QSiJUeIFM5Bv8b8h5g+AFJG9+TX0qu1vtow074J/2RGilGrXCxAgTv
nBVb+OOGCFtgM3NE6l+oy7Pm+yTFMx8gSaq8WDZLr3cycAiVfAtxDSahk90kEXZLqIZBrxdOWl3q
kEqGuD8qCc67fnd3TQh8c5pYQ1vaer+Rsc60dck2ayDVjAnSjS9VplpeXwSeaW6gsGrpcgF2l5Vd
RfVAjcN6WroZkJtdWABrXgWUWySZroRzssjNq8qrQL9+PmF7iKi23z9tbm1jzZJMJWPbvfQiKAOZ
7719Fuz3QYoj0dVOaVlgmSTbq2O1LYsP6eplee99jhy7NWIg9z9UwGmE8hrStx+4ckRc0z0XoYQw
Xe9o+JVAG63+6b2XGxEakhFxvP6QmNfbkawgpfiBarsWSYp64yUmr2Jq4Zpb+iyBDIEHNiwHDta7
Be1vB5Ot3Ej0PY2r/u/dj6vOHwuOcpKLgRXEneEcKm+1Y9kwX/piHSVbfN69rH6wKx/Uhl2pNAtl
nq7cOYUj9YNJiuj+ZOXfqIiwN72cte02gi5OmVN9lDdWbdrPQ0aeq/teiK/lrXXsEB3VzKrWAnY9
5qT63LFKJ6kaQzE2hML32P4vtlELYko8gC40080gHwlSmgaeSPLxXBgXSAQRuPYh4iiDvmxqamI5
Z66cgbr5LUWW/SCEAYX/pkirSk0yt9jhuTpJQesS7a/EhJBhZ9FXro36qc1KtYYxakszX4DhMESe
cGY/oJ89cN7rcFXhpiPjafNyrNwaDRtz9i9Fhon6s0weh0RgEPrtz2sI/TNzJpUrQhBJV79uDoL8
ftj0TugzoZzj5iOyebtr/sJyT0nkmyvsTvnWu741Dn+nf4n5+vZ/Q+4dhJVfbcaf1+Pi7d0/21ZF
hXeFoJ34dfk8KhidMnykF5qebpFG0mQoHTkndn/WbLVZ9Iv04yJml1HNksXazLKxf1TCi6JUmSfW
he396GFNRIoF4N3gsnPpGkOKQZLRmoRH72tMpI8orNwxgr8Z24BxYhTacYwNnS+mRekl2nxguiNr
Nb37pwRQFSZOoa8dZz5z+FYIUZAIU4qF2FpGZvwzIaXVEQjpTv19NSLYRSbX0To4n2ezdYDGziDF
dNXTW6f5qJQgG1bwBebyIc0pma9bsJM3HF4wXizZvo1MWl4GBia8DP0ty/o+SUgsdXfnh+42G9T/
uhczrAJ7oe0hGaxCkAytrIKwv4krfagAywE3SXDlOcSfjFA6/3RN7DhVZ8CtJHdkjH30w+SJg0+p
ydwWY2VU+7mwy+amWjb++nqy2P2tektIb6F3mfWcaHHbK/wzHh9hwTLB7E2+toFKAB3EBnmhvDGp
qN3B7KLUWTLvmZV/sPudAqP7V9dYFfUy6EjUE0VTW+NJ+tIAe5VMrMzL+guIK8Yozf3ks90bkufi
JcO6oC37ekAsBuZXYGHSvS8hkfPxOEy0d4or/fz8jxvEePjBb/ZEjUZdM4NQOAtyhrceToGwto6m
Sh8YzYa/dcr54zu1dOac2mj0vDEeFl+KqUPYKvWdjtVgD+aUBx52rQbHX+8LzfO+ZHa75ZRPlUzW
zOW88KcZ+qEMopAhcZQipfoxZTs0uoUFep15ex/L9ZhFNG2Pxp9uRNj/yp29cwWX5XA26OVAnjSf
3q3Kk1SR5QoI77RO4AbiSDBMCgdwdm4lneMgrDn1lXJZfiaQKqse9ihAJot/EknDhPrNEv1dcfEC
tYgsLIpRf94FMTfBoqPZHnOkNEYbmuBL6pBiRC3slf7byPg9O9K0cBR3XMmmjoVju2bYDhB13OcW
0JZOOMD6htIKYCtw1Bt4XZ8H9gKkFM6/5/spLpDcneAhyJTY+QEuRgnOKxLRcd8C+rwJEErqO4+l
VTo7NpPbYhGOLUjU8i0pNiMCRmDzVHiH1ci7jSn6xJyE9wGQDf91Gl8cOQzk2E4K5i2CNo2WDcLh
Cqn3kXhAuSJ6gMjxCgvI3wVozD1gUV9EpumTZ4KbqnR3GHgWNfC264khHE4vqXdFbMDZWqwlLF0u
xefe5gqav4l3KT5qP4S05nzFUkwEhFUSvjL/AecAMzAnzeOO87scTK1+aZ60sz38sDL+BSfNc2BD
IwHomdmJpIy2bbafMAp0fasIsPLlheZgMZj4r+JT5f9pqM2QFm2q47fd6CQE4OJ/u069g/p7pb5S
IY3scEn8HpcvU5FEeB/l2j/ske1wAzJMwXkQtsZArKHeZj6+T1BtkaOr9YrxbuukvkmJYktNh2MD
p0EjJTgp0Ins5g+oXJb34m0rSreYQeT+1QSsl5SEBBeEUIpJCLLq41NAPhhceeHL3Q1MZwMT3nqs
M1wzBIRo/jA0use6RM0yUGGzGLWXiO1kOolUW+idl9QoW9YtlCnZBUoz+Xr9JpHXZlqhXh6TLQaJ
f7fTVLeXayUwSWM7eaYXIjYzO1429MP+SQhc+haKroIlpUVzG4DtpK4Lsvxkrl8KxWR38l8ZhEuC
bRMYXPh1ySdJUL1Mx+0a+ubPZPMK6jiL54jq+eYY/LF2oUM6UMPGQyWY3h/wQ+oPNjVpNLrmhjFa
IcsMYTECkS9/gW9wSn8ta8pqeS7ptNWJ9n5blXK3CSo4+ViwLuxizA1y2DOzu2qFDB7TOoseAiIG
JNPsnkBInfXedbctUmhoQW6kMGwDNkMDGeoWSdjbGwFfeppTyuJynpQ4r6FuOt+kBUf/2HO+16qf
HC0ryjYXDClh2UMpr1Z6qOMIDCKh/1Z/q2ByMJGERl2adlkvQBrP5nXqZpRs+C2nbbBKUGmedP8b
jiopKFG2R2EvC2zhVBz48fJxhNOzWuGwywtIFbsCl0C5f+QOaAlbh7vBvsU7aN/KI1g5PAz/6Svb
CzSsJUwQybpu7NLzy1aDMdzt5AQ9BWMHloFpJ32XXOBNfqPJWfOooz5V5cM3tF3pqeRAp1UHA3+D
h93vdxFmbfWs1M5VBqUUYFGdzpHDgj4NM2uoI8Ri+OGh+ohG28B4kIfhiRe/YwvNKIC6MiT/f6L5
rX2wGKgMjVqQnnRlPBfWdntuV4ds3aE+a4/8BaTz2Dsk5eEpS+9g+CyKPdue1v7X9evJB5X9+N43
h8lcRrBuf9IFKCK5khvvFZAzqxKkMiPIg5s9vdKS5w6XV0efN3X9wLTZSjOOVWGtQ8ruiNhsq65D
OqsrELbBJSo3aMFfINTviOFx/n6WJNwCrab5/Ehvb04m6piQpVnmB1mC27rkRxUzHLeg9s5In7QI
cl5N1MAC3HpDyI2LeTog5TusGJdlfMqeQ7ELrhs18iSM00DcMJ7/hpVp9wtwoZzjbcFK9CJqko+f
QyJAas1Ng/mndcTj7ucShmjX9HpizmTA7Fr8XG/xCz8NZeIYOJUXAYSPIjqfCYDH5GzjXMx+hAFM
2mqF7bo3Qg9EjSsOoGpC/neMQNwjBnv80tbfPJkicyq1cJ5Rq6eFwsbpS0FctKbiimubGnJ8hmWt
K5ETmWr/8tsi3l5kPl7FwBZDXvHrA4ONSsSM8qlIKG0+axpipg/dk5oKIbyD6Bp3Lp9CSurV95Iq
tSYeGKsYvB3N50z2Zs/uquztMnLnTRtQ5AMrVHZjtDgJ49hQoDrEDtlQIx2aZuEVYYwFTwtOSkjQ
1OBfPAHNOWbmDf+Mhj5DRzWSatqC6bRp+66kNQyH0JBEHO/lBgNzdnGmx3O3rOA1PoKqlqUkgfno
Tjq6jS5UFo1XdHzPOTYJF84qvAWZWltj8i3SPCJdPXTpZ1LKU1mBrU6Np2PpezFG92QOOGKriTfi
6oQUa0YYUA0Xn7YGa8I6zrKpeC120mGZDPquz664mN4mMXsvlH6zw2/qRJVfelvARWW7VFniym9G
/bQCky8qrtk7pBLO04X2L6ueFd4S6JXlWE8A6ANnu7Tpc6PYjey53dVqUKNNhaN1HB/aC5ZyjmFn
D1v1QQX6fLb6GxRJK7AiIZnayPbhRc9CQ4rF4a850A/hpkO1OJv1f2P1gjOcdYKPoGAe4ZnDtowW
Bs6h9rXCQRUvFO28K7bLjkaGnLAPEriEqMt2qsJLHEVRuC1Gk7cmFSGX6h+0TYfYJWRnOFF7fDDm
KGPwhY1Cg6NZfuqA7ZavhyIAmb+Evep3sRwpJCGJevawc5UuDewHQ/CHtNXabnU4rKGWFMuCZRb7
eD4Lle/ZM4EjeZ8W/x1+w1Fz8q6h90QmfCWELMy5jCWJ9sMmfBzNaLppC4yu6i7ep8qnXwja/p78
R1UtQ0QrLapsZ+0el9/X7MnM4DAJmKrdwBz40A++qlt3t8bvdgZTyklvNGDf08W+c0rbhTvubTEP
xH3gPNLEVeX/b7x06agwv0Ytvh56QAIO3UjuMl3QDky+HD4ArMCWEyiBa5utDZaK25RoREEi6wuh
QEhfFeY02AUb9qw8OEhTyA/nkdcg4iLnv6ec1w4ElLdA0BrmhIKmm49pbci6pPtYXyvaHoKLKmG5
YvSwVfaY0JIti9fYfxlWKQ7vd7vcBd8M2D+2smfNrK8hxb7ho0IwKgDEmyBIiT/6FRqWAtk/XVku
IacoJp7nEBzjnwEbj2+Iwv4TVBvARiQ0XljrZrmMWPDG94Az/DyjPsGxB8lD+bKlSys1xI9ijnFX
JbWeqz86HYW744OXbwpJdvos7AISEQjM86VtaBGeF5MX7BWAoP/679TfymKXamHnUQEXV/tHUFpd
htszzoFpyy1Jh9rGO2ZQsjhLDkLy88VJjde+Zb91VzUvpaBtJYlsI5rGHm3lwEhA5MUPME7jWtix
qDG5H/i9IlTWti72qRv4CiRhEWuYHwbYFJnwT3t4f/IdEuMx3mpNSEVMOgAlj+7/wvCX7yqGZgYs
wNqawUaK1gCmlqnbrgDzmODy0CLA369lCmOpqNSZdVqxyn+AybUnggwNdTz063q9ExKdQ1IqmZyp
fNU8ZKq2CYW2CiGPyPvVk1+RC74HB18vvCwoOlCAtSHHgT+wxImr6SkvOhbjM8qAYM7SLDbU2oAW
6QVZGCKSOW7d9IMABnnth+PRhd+UaRvYaOVqjH5VqUlIIEd/jWW3ZyBOtlo1uiFsQjyhNouzWv+w
bbxISoPhCKWxan2vxsrLbjDutwLoUhfxBZbJu0PquzpS25a6oMqBp27ek8b2zoWlHQfHwk3AubRz
agU4zJe41ipFe81N7tTlmyUy6mbzYR0FceIGt2QmbzI8iRyqD8aRVPgrlqH5Md6S5icKPlWN9UDa
qBtDh0oHj5Ae4cauIklJzNmRbtAotsH5CCpw0Nilhxe60P745MFYOShj9725VIRfwDV6tEWX96F3
dzcwBNjVb5kKPH31FwMYPionUXUuIiELBKUQ5Ka5ttIivr7o/jOG0um5CT+RBH48U73DBaQPR6dc
SWyxGKdOkqO4IflpqBrut7ESAssAb3m+z9GzFhfJsa3uO2+Ic2wxkK+e/bOBMwyVpqPr16XEeagg
qOHfYOodJLEr9JDDHG1FdoGzHK/CtfypfU2mgtxzAHNfQtoYljLDPWiP4S2hL01KbkTY3k/hB1at
i6mWhIptPKuG/9uLzb9iS3hBUaZgzieZeBVCaQsoPaIJ0g/V8om70lyfyVVgO5ADPFKsZRRUg5x0
1pzRGXQc/StKDOlTPzjocpNunlLsuve/KDIK/KOaQYcS/m+jiILXH/h0qym6iAP5B/Wdmwg5rxDo
MPGtoVvaEe8z1O6hYicTDVAPe9e5rA+SZo9YoJini9sBpgLwaTuKK2teUlu64rZEMky3X3ES3hTo
9C24dz53G6jBNI94zJecfu7Tc5kgFpQb1qBJRnM/Ahj2MZvyAsfVBCIhYg4IPwoa+961W1Ih37Uz
7PdQaHNAo/qVZHPHVHD+tJze/lfgPSFLcNW/LjadIPyPcLA7XILuuG04X4HHMvSEtLi9hgpukuCw
Y5gAMbUxkf/WgOi/EwtquDqEN+2yK5vx4d4SKNeQ8/Db5ldNHxJKw0nskjcMRg33eS7VISprXeet
3Tv0qXzY7qB8LcOLPvWpM0DsZbAvO18A+4nMv2HYvX/XXoG4RcvDyBVozGisYZqSL7GmNnmVUvLg
DLxf7Zcq3OqpP2fBfp1+Qz+yNXt8rf2qwg9DGIns128z5dZhgIbXSKWG0+IFrO3rr42ijUsLek0m
KdBnM9pEI1FHJusru7g8Dvfg7JMvbV/PrqjKEEhZ3I2grsx7ilkN+kHWjc+Rin6kNFOS8l0MVofQ
Bumvp2cx/SzyD+tte//HfQz3LmjK/czQ6gxHBFq6/eoyDzvuxB+S80YidXGA1Ym4IG6xWeQ6Aa5a
YyYY24RH/3r2ysNu96LUpdfz4+kTiD0+H6eL5KHvmTJ27ki8BZorpwFlnQcDHG5xC0ODNAr5dQQk
WwOhV/sE8ib0vinFJQ1FoSXkFlf9h/eu4jmOmfnJm+yEK0EB0xncsEw96r3lNwmJtav2a7pYP8D1
g5R+u68HjaM7pKvUoPb8EOda5ZkMdwGou1z7f3jZ05RCSBpqW6HiXGeyj2jF5zxQeW/1xfkgmLg5
2TPKKNUcK3l5+uBAWW/G+qClFT8Cmltq3P/Kx675EI8JRz7Hcz5faoVxvR7YO357MOvPt6uQ/lgu
5jQp0jAgQnKDvDdeCEi0StGI/B/bY1z3dtw1W2aBCol20IA4zgi9ANaS73knpGVI3GgltKhIEJug
LbS2qEtBXVxqwECUB0go3b7nDJmJNOMxiMlsFeGHEGwzyOkzL6XsknXCmNmN5v4PUPuOBHTYVq3w
m2fuXWuHuYbRJMxGCDkFs+WfrQbrvjpITGHHgA2icB53OyUGmTJunvLYcUD+w6uqL4elWkRFGMke
fa6IYQlaqOk2w7dhZpp83xZWSmA08HO6D5BIIxGOtiwWwZxun6XJlask0wvJfN04BPHQAurGV+sL
uIowfTz5AQkm0nEf8mWJLsCQl6GsN4oCdkN+Jf8tNNKnloSM8pmx6g10qgSFD1gjxkne2maOH1z5
zeAIbecFEXp8EYLR54LDd4rcUyuMQ2ocXjibsr+UgdLWO9s/dyysClQx1NDhDm9G1bmHzxN0RwsK
xz8mdWbFCdWBc5by0zgCMEepq/X4p3UfDK97/K63je8KzhmBYuzamWmphY1T1aGHfFwbnzNWTY4z
aboyjZvMlNBLQUe/3/T6Iwx7AGQS8F44mRxjGt3gfmLqaKkqcNhdXu4nVZRqTtjEHVQ/qc5s3VJf
sJXsoKdrqdoXnSU4yxLrLSpOGZgJATD+0Ir5X8Rc11L642s2QGXUQH3oUrx7wM9z9tBZezCUbqFf
9FCWNFhZ2ldb1nQQRm3mkFNXWoM4R0KNcrDN3QfSjsJ4DHFZiz1r6gxuYS4rbDNxaC2YHMrcXymp
uwJHqw819M7kryBqeymW9u0J9sU+6Wk2aik6cEsKWdQKhxTPsrKDIoGEvl28TuDhyj3VLODbOwas
reSC6xVx0HFUA6VtruygpdYeN77+oxcoj3rie0KsERZIUJUe8nl/b2TqWt+Qojq5aXe2qU4wSufe
LX5HxzobeenxkoAA0sTTcCuz37bsbzYSCYIa8gntg3ds7ftzCXIdQ7UpUEpacp5wesjcYgvenLUm
jmq6WRfCc9iLG2KoYP2PKSq7Y/f8xEPfIIw6hO9b84Ga5rQF/k3/e6wWEpL3qNUDdpdCs9AGzXLf
3MHrPZAQR+oomfCgJDnC/OxTomFZf0UDkxwZuK7me8xZVaskfe03GdpAqlW45G91uhmUlsT7fA2S
WeOgxoBa6DgwhEKFy/nJUcthX6ZmoY35Qro/iRQ5vMa5JQSta/Q2+Tz4VRyNrINmAcgIE4A21fXF
w1qZUcbtaQBf2khprNXuJdEcYYGwc7PSKfP5EKWQ4uqReYYkORaRrV4hC+wTZR6ZzPk9MPdpbs+u
c9MsT6FYC5gKeaNOK6f0gOnyAFlnBtp31zijKpLKMIwYNcSsqxGT/bxBAhKVs6PE6ZPzglD6Mu08
n/lclwKWMUO+XTp2c6lCnK9fJ2OMzFbVtcNkMyvW6NDro6WtnpAnnOSKqX61loMrshZtMetUgpCB
wSMhOvvD6x9tdgmo9oGrvbaL362JSXgggpWugM/Wqb0NEfMvGoU2l8Spl5J+sFFz5WVZMUqx2hMu
Di/gRnI221EpWZ4RO1MnYjKalVuDkri75NsSUo715LRDFLP13n0cbj3b9JF3Ylv4mHm+OLvNQo8r
kNElr+DS+U/6OImsQCjdfLzAeWuFFEgqpEl4M9JoMDryabKwi0pgt8f9EQp2QGZTIbdg3QNqF7+V
Rkw2O6xUcHFzoga+eIr+Dj2quAtj7mnveQhJj7CF1gfQsdijmY9iR1Jq3hDPm8iMkFRj/EbOdhs8
O2s4pQpojG946oYpkWiWoyaIsGJgHks4QdZA/yXA4MQVNWUgNDW8B/21yv6v0Qm+lZksf6fU2eMy
PW6/X0kJmJHmK++1Ii5vms1rltTpHWvJtlzadcSmHzajA/DbBJ+WwQ6gyq2JTgfy4P5ByU73Wpd8
iGwdSRMO3JG4Mtt4Md0JZmLzZyjfuBzzD5q+/5WlWYtBNE/ABupgg+CZ1hJ6nI0WDFa5UqT7796L
izC5N/6pDDz5adTP7IHvnisJfl8LEmugxdgLoYqNHW5rrE9ySelZ2Tnr+Mmev/a719IRMStYiMrY
w+xn9wxnlg0Bh6flewqhJngWwI41HfCoemAw03ohmo4ios+MOIlzDfEz+aF42ul460aWJiIDr8sQ
xLjWqRtn0M65QVzw8zKGmqm+SAzoW8A6C9tPz1XRjkvLVWLLs+gdgaZAm2sd8fH8q8X9iVLmoWI7
V8JS1PJR1fGt/XjeTKpaA47VDsH6ZtKKH0VtQFKwXguGhHNbbpwE6jPHLPQ6M/bkbdpx0njAzev4
cjy8W5jHEE222b1KgJUXHToEznQJQf0/B3qE0JKAVJhA4LbXcccN0J1h2lfMRMZoDPEDKZk6aaKP
dIaIB62pVyTPUE2rNxwuscHgqg68xPqwz6DhgC+UtYZG8WiPomIuhr9BXXS3mYmqOSlvzuvW7FOI
RFGTMr1xQqWUqhjmLYvbMuHwCHXgfyNMmTkf2ptgcUHQO8NdiBo6xixy70HkM4UPjHyRj8Rcp9XY
8mGRX+t6KcwIZ5O7Q6Pbx9yiePmf3AtfQwb1yQEfKF341fRa5mtCDLwZeBwDmKpHDdxmZTj48vQ+
7TGXFcxskFLJKPT4iuwn1I00IqghR08cA81/Ot6DnexSHF+tVrWyC0FeisEL2EP1XTArhF5/BZDL
AmDtJDdBkYk+Tj+3RYWgslCERBkLcYs0qOh0+O0+qQmIr3rXiogJiBr0T8RWPnwd16JnrJ4MqEe8
0b2QnaHQotaMSvyIl5NcgBDhi+dHxPjTWYcCx+qv93KFgsYT4QQTlrMxnB9g/bvvsWkbCziuLy5I
WcOF4foXPjdGeJjTCY2Js/TpclCPKuIzmIIGRUQd7X4Fx3ecrcBjRYwqKtvncn8OzHgemx4NJQt7
OylbOQBs4RiWvcB3zLNk3ksckahY638KC+ySvDVeq//m+nXTWwWzzkycInbIiHYkDYgnbJalRu/Q
+go6HJ46W+rLJR4KUqud1DKoFAf1DX+URKyxbl+RWRd7paEInoSGC9GldMKdzhrKGumckIkjNqop
cex+UctCUWOLXbLCkyey82fksf3sCU4iKT49g/BAelr6RCmUnGjG2ydD9b3iSRihhn3VYCwI6eZx
73AzbI6kQBReWAa6jWgiyD+0sUZqZA7cmw1prw0P/KVqD0FP+zs197mB3D75XvUOYztWEm8FVYVk
f7Rk6zmYy+3ZoRyZ+uBV0C73YH8xXGlQX9y1BPO9rGQKzXSPJollMa5eil5XGo44zDms1rpYJaqR
WF+xb410EN7jV5tM0v7hLRfPuQB5RKXLGLcY9Gb5B64OaenvRJSOmunp5m31RRvvL8rBLeB+bkLC
YFQRgNKWzS6OKXcyqfhPZYYs6fug9XpY8mZ3vYFPRJNn0TUoOA5aiqZobJHIAizzMosr+JSDdTAP
FW1nM1vnpxGQsdHhWD68SZ4PDWEbNmdp7QusT5cXFFznx/olyU1Vij+6wc3HRd89uFAP6vYRFeCm
cz/+l0+Ol29K4O77Xs6KcUCr0W0JEl4vm2oaJfz6/usEvJ3RGraFlMHCsX94KA/7WwPX9HauQRPD
yhZ47x0G3N7J3OMzzpPNBPLMFZv3ONrjto4v//tNjgOcLJfbexZdKU2qCuGdiq++kwFVBL7LMlVB
6cno7Kje57GflHgE/Dd7Emagp7dktxXqBRdALIXA02wFuJb3NDTpGfZXDdRp/7rapl8OwScF4eqS
texFWUu9sofH/kxqKqDKBOs7ZgU6BdNtTzOB1P0VdFCJKLaU7TUGUeaQLzabnoG7MIHpqcANWq/a
SqZNCH7ZkzJAO1+O0X09r1dyCIF6KiONmd3uJPW79AzILBULtdqY4yPVxTeNKB9i1s+NT9LYuiX2
zw5+jPIowhDoVidTL6NXnvMTeIozs4g+BqiDb9wb35wmCrlQAJ1tx1YGUO0gVK2qv0lGMkqV/Rzv
v21aVjJ9x3CZyer5przNvPNNNgWll2N2HLUIGL9afqET/ISbkXehCiT6XyCOlnxuZjUdr0y4JRls
L4R1tjAIFJ02kSIoCyad8+WzgoUGl/yhHhe/UYndiO5JdZjHn/Mk0gWbQR+dRCpaLataYdG71sBB
2O0PoSLAlamcmt76t/Wz5zu/5OGPIHpVChnFXDxTVwm8sGpU6EpM97hUwUJHJ58otIAoK3fOjnUu
NXoY7KKqtYyTRzqP/qxPsqEqsfLU5n7/Hl5n//jwHm9NgEDSamvrikpVOI4LoOqIuMtI9bFNURKA
ey4W/R99hK7wEOuV5xWMKgWLH8QTnuVdpohjSbp96+xjmFtgoh5kWrLC1SywT5cSfeFfqQh7ZYe1
tLWUwmh29YIgIyZCjIyFi5JtUNH6WCKYZ1hnQJCkQ2me4kmz/P5BUSoN6UzNxisXO7SCv4rzntHo
VqlKYLHA9xytksxxtSWCGJRmVCRuE+oNXGx2U9LGz1RdfSAfcKg/MBsKmYQZOQUycbt0cyTR0pVU
rhVZm1z/OFJ5AG8WFZEaE7D0Iba2HNgDKq4eWbElwCTVshtzJ81zfGxM16DLKOs1gu9wLtYWUP32
NEXsLB4VMnR0/g3T6A0jKHoHplanNn/blvQ51MQpSbh8kYghOZ/S5R8cqMvhI2ADb5Ihr3k1slTf
oJV9FQUQ0zeze0ikWBVjjK2n41qeGp0NPexrwW95NhFh0RzDniNiGFPmzUj3nFahKr4GZ90zeJjj
e24dFeKZiLZ+cyLggQpRm2l0111usKtyzLss0wvhyOykdvx76M1QSQd5KCD/VBpjbH28MibsCVM0
JHmjJBmqUcHeRkGeqsAtYsOZBXkR28o0QLgkQOWNH9qQp7IAezjjtVzrfTHYfrLWxoJtuUS6xaxp
x9ALaI4uNKe2M9UExMMO9A8azK46mTYRg5ILUFLpMgnjBzJ/UkbrP0e9H83/mki01Trmn00Mc/bn
asz1lsOInAYyIMaDOura6EI1OkaaTimd59vGQoHWy4orFWXJjZGzpn3KmcRebfMHZZtFPr9z4cxQ
mRp9wUtQsWvXezzusloBGj6TuO+nIgrX5UQ8RxhB6MSIouxihuKOBXBWzDaRI4iU8yW3a0oqqEHz
rsdv3hMLhOt43+4qXeQJz0QI5d75svOuSCOV+sIIZ4KHoNPnnw7I8EDb7wEG0inPjUlLz6xwG0yG
ZfhGamg4WT9VRG6c789LQJX2FYhzzoW+SUwGGCC+xaHsEUPnIUv7WR999xMP00VOLo8sjjki99lB
l5OuNQZEvt2PnjHh/QzsucwIx6rViiBNMvNXOUBwsQbyLQqxVEAkCTSoCWiYHlyuQKAVa7ubahO0
DDmr6rDcgZGaUoMA1LHnUVp4VkCPMJOMTEuFkemn7AOzAdAiqgilGQh/7N9IJRojokYqxyYWczJL
gxwtrVpkqDb2GN00QcnjzxmwGo65PXu8AEHNnVGlGemtZ8dxMyWmCvUMlLDYHdWzL3lnwpyiNc2u
jejs2QJY0OOgMJisVqzVfc9L1F31yLggMPIsjO41Vb4M43wp6vF2mjRrM6fXFEH++uzJPdsrIj2O
siZjqqxrZitadJTwaUVnjVc4ISG7ZyZMjCMMRCctuVouqATY8r6f+7K0RUGGc/8vy57r8fXCauSK
fXh3AmzbPe+sdRPZ1BDZ6mkrpS2tkyH+Fg3ga+Rat9J6ss8NOOlwd7mCSwAu83NE6p32y9Ah2aGa
19W1fS0xC6hZJoCoI+w8L+uWwTt6FzjMOWEl9iqJoDJ1ifqWpq8wqIrh5eTeh/HGebgM415D61PT
QAgzCSPc3Silr0E4uGcFjKWoWLY14osav80JVUDJJDzrjDg3OCzpsavpv8+yMb/S9Ws5BIjuCvPN
p5oAw8Wt0OPX1NCjiDscJpk9CnQFN6u4KVeqsDLNrUNFoE+cYx9Rf+jBxc5zxjPmGanNr4DzhLzf
eVOMROrNXDqmjfrEXdgtClaBPvAyakE2D000K9pI5TVD8AhgEzxFPskAjVBIg7QV8QErfuTVzAqp
CN/I6E+JZnjy7fQGTczxSkPCeSWirjWcOK9WYoQJA6GIkzMA4avkMRMabMcsc2yg0UDzlPXqvuZC
jm/KC0GTV1wSM1/qPw8cslchCGtiz3i5oe+GNZzTpL5JevFh+ZYvvyQqCpksAGtYm6XqtC1EZ+SU
IudOGgjML8swzlfPO1jgS+hPBmK23mwUYO+NNFIgobr+lWX/FwS3Xt0mPFtn0GZ6k19ZARxW2xBj
BF0o+AdoYFNCQbewEUrNvSI+WQUeGmwv1ahUEtir1RS5R5ZI609fnTiOZLTbjHDWmOkoDLCkNuyb
tiY711otg+++IORY30L7AykHsl8+lsunE+PECV0PUFrF+qef8gL9dtoJ8XfSNodDcvvputTc47Wm
We9lNn1MbAZCfkciSqC8q1Y76tWhQUepOG78tXTJSNNtnzK6DcV0zYDSojT7DaN9AbGUCizn9edy
PllGb3hVnsY5c2dCPZEUgD4TVf4mr+9qJPiZNV/0jJPWFCzkRrTavzD70s+8RWxfmoKg/WSqIiTx
ojJeDKDyGnM4a43pcwZnuRic7gQ0d+6R9R3fw3YYtApX9NmUB1TEzywE/ME+foA+ZkMX4wvpIS/G
QUerQxXKqYt3x4P6OWYNYxcgPkCqBkkLQvfOl9xGCKPvDlCBPISUMIK9CgV7jSsrymPl8eOkxN9A
o5YCRz3SXh+caALR1MOuqJNhhYL7BZ9CkroULcm4ivdcoG9tyDt+vtQjPBO9khPuXoMHdfpVnvgB
ZrEhBfvuzelV4mAIJtdzdFyJWmrZ3cYZXihzLAUfPwvItxn1PzQ3ibgnPwAo1n5tjGExIxUKPO6e
YndHB+x36x/w/3IKu4twFJre+Iq7WXVXWDLYGM2cQ272hojVPeeK0YPP75ljWn6nt1LuNhNqL6cx
pOtOSOgasUaI/cblY/VM3ShnT9hPm4Vcv49Xv7hBylLTMGrEAJcOb+aNyGfKxKOliCN6BEIofchH
tOFCp4MQx2+LPePWkX1zYJFGEmg5JuBQYQxUAuHnvpGPXuUp4JG7N4slmf3F3CW8gt/Siv8hfa6C
2AjYkPJB1Eo1D7r43xOHaHEbgy7ktdtiypheHlP5VggEi7v4YwgDqHdkhy/3gmyntqowvGI1pI1f
hrBiSovKPIekTlMGxkB8ZISJvW0+vyfbuj/reu4g9nXTRntJc7XLVKwRvw6jWUMS1F1Ojgld7Mbv
ZH9a694HQ+AfZPZ7PIjG30ElIZ+ZFQ0j9JrOhB/P9BKGacw29Oe4Si2otHUPoDHCpdZL26vnQb9u
Rgd5n7XGTKeM2iIl006YojD+nlt1P+pxRgdZF0bFOjjv1p07/SlUkbi4mFy2iB+/vA+E/5pTHOSu
RPDNTSSiePiYRvC1v7Z67Zzb2Ab3C1/ksGlwD2u8UNsBdlNNrxjqEYN8EJpJLpdQKwAATYIFaW5b
gM3x5MwAkgPZTMM4jvhTtaKxQpom/LdL+K3E57kNABYnkJm2eyEDKHxILoaBOgwWbes02Tz1as+O
WgjpR+a9sCsKdmiD2uDC/YyHO+m+c+QEmOOAzOCi55YOl0NqMdfHvj0qzmwGSK9S+IHC/zR3W8dW
y8BjJ1qdVfHyhlt8NcAQzKVsGA3u2P6G5FnS0oJtAzVMpfbEJYnSNcwUMcF1QHJiUEvGDOY6Ts4N
pj/89RfnCQrwPpAAJKM3LtgBixWKeW2j/eN5AMteLoRyxWK3h1aMj06BijqB4L3AV1tGVx1Nzcz6
wR+OCsR5/nyf2PlIy9gL3X7cpTyHz8s8UptUyJhpvYz7QEMYo729RvjWkMqc0AFK6s/DafM7yx5K
38rQa0t6AqMiWn0DBn1fMyf7H8hBQscg+zEpFNZPDzc5VkamUBqbvjPG8Ubu8cdIEQEci80LmEcc
UvreRss9Hjy29RTy4i8MFs7uqcxhafnHzJh1p1RYoQAuKBfgMmE3vaJT3AeCuBukjUWIfa9uZg9l
PrhVJ8pqAgOo08dxhxsXa8FqpHpqB1vvl6uusEezt08VT6L5unp5cr99BZs+LMHCR3x/nh9frC/5
3RtzbwoxAjyrwVErVNycfIutowxKh6q/EBcULgL1lpTjE0WrKMV0ZCc8VninXZdPU0EhtXFXqhJr
hC9tvktcxzWUbth9B5I+0vWpxPFNcWe959ki68e3DpWrCN5vHnujGdGW9i4mGSFJQe4c726qZcgB
VlLvdZPR5BsJJ4NDP0SNlKeQQ33e8Xq20rrWKcSfviyZsbvwtvOTyHFUZhb5fQUZ5vNTndlqxNfu
9ZTkoq5ISd9YqLa6pyljCMLmEJW9b4ug7r0hEj+pN8PaFqvXBjbWu2tiqpzeTTIXAoreouqnNa0F
tqDd1KrAMeQTP1yUykaeJ8CfNwav9eUf6t6OYop+GGMxSyGNSLOlxdL6GlqkVBoo0HHDIhatKruc
kJKFyWA+X6gM/SPWJULFl6uJWhNLQdrRS6LB6TPYq4lACjkGfJSrsZdcMM+4PLN8Zf7V3JnkHM4v
aDqOnkk8XnWrZHKIvRWjncwE67X3JPZmEI3JrpzncoLju9JbirrYET3ewXBKQryhn8uPeuizPGO1
h+4XvSWLHsRx/W1pv5cdrnuOM1IDGZiKdq6vp8CgQxIaYINYYg7pxeP0l15uQ3PhKGkx0c6773IA
Isr0qAqhzaXoELt9Vpv/51mrxgfiExZ3Mvl+68g5gesBHsxle7GMuOWgbBXrbnO12jnQmAClt9NG
4klIisClSdgOfU4bbwPi/7dd7jRVIrlEwhZfDnQsWOxr5jMSBV0B+073JvKE616UJmmJPNOLKWBb
QHkltq9ha1PfEQzzbzW6LZOFW3xyqdRZnY6PdRlQ2G5w914/NKvC1fHmYcpB0R6SclAcKburuEmS
DbZV8PcPeEypgjwtgRgBcedFEbBfk+h6RjyF7AqQqkAmWgkKB/EjNCu8WXqtl+cgWf91Yq499uHw
RVHY6o1oqkcScno62u9CqXVhRCEKfqSgJNUk5xSefW3BgrgfYKmNHrHXLapSLJN0XEin/bvXDulc
5Ulu8OjWJCPklni974hwVZx/cIZTgTyuqVVvyLlzfNSDStvvOfI3DRimxeUkv+H4M+yh0jYbKZiw
cvHyvoIGJBov/6MbY6uWj5L4XiwfNgH0TV4d8LgXxy7a38p4co2P4Qwop0EQeh4PB1zmtVJBQGTj
at3fpIqN562WHv/EqilM1IyNVaKnzEu2v+wIG3t/8H9D4DDR+xs1W9k/mcSKkF29RABGRrXcykrP
60ldohiAgdlA0VlajdRvDp1zsqLUnqkZLg5zUrEuQRgBg+KgSbmTsy98f7YvqBWqWXMClwtw5c2X
TohXWZTK7MP5e69JVgY1va7f1eCFxMAGHddr5vzC/wqNgsG3ljjv/H4Cir6m/i7uSJ6oUMvbsEaQ
LDAkjy5EDrS46jqsKAWj+7pZ1nn+sPb0oA96T1MDVIPKwGiHgt1JeuzXEhch+m30gwpeeGlhwLDG
LYgS+ezAA0mDGA0S0Ef1hpvJrtOdTSQ1hhHcPL1NREc7hB3c6nY/MX+dHnd8LG79KsNpLVCgtKWx
7+jVNiKoCAPTumXyENdrR8KAeGakVtOicCNo6ytBcXCtJKA3AbC9oMe4OFEVHtm4uOy+hmFYhxMO
6AHibyq6Bfw/DYONc0+W7TPR4jb2t82/1nLiIpfXvUsbqhARcahrLObKxCTw+kRR/o0O21PwGD24
wIOfmIckiju6mgBI9oWI0bWyvz0ymKJoo102vB9oeLx4ykbcjloIO516tsmgTET1kj8gLlFxN5TG
itLnabV3+E3AJzj1462xmcDMiHOJXphh/Gv4C0KWMuEZy2L1QUm6t37N6HQKAdQi5/HxvnuGo/dP
8547IzTNWyDZee1QEkFx7QARwmC5SAzn2xxLNGj0HBXmkHAviiwwgnISUa/0UH5GSP8C5OIQ3Etd
d1E0qZLU6Iy4nVEF2jIEUqHoc4Ef9IzJNEDXTzwb33sznkaRKi1pAsQcE4EMKffa0KoKWpiucVeh
CFv2UFyt+mRHlkWLm/KvVbojXdRQWBdDLsCukTllnMPvLB/fBX0zCsD+9FFsX935hKs1E2VGy2sf
YLPOFr/qSqMl9eGB+hYcMo5XmwywGjQm9cEylrmgu0l2SkNgkEd6OT++RKnwfiuZqTT5+msa1bhF
rs5q2PFXoDJufwbkajNLRbZLP3ZKmiU2JuTyksBQyjlnOIymdU58VYX9Ulvi03ZuT+Zt28RL+Yrv
b66cqWxHZZxCXy+GGo8/OBFcjcPON29iA93BhDIdaXdqpdPxznb+/+AtUFjwG0kzdVI2hmr9hDqT
etgWXGbbinaX5Izz3l6zaKTq1Ut6h+2b+1mDCMifQkmpDDg6mqfuDzd32KC34jVoRZEi7fFGl/PZ
jgMZjRPo+ePnMU2l2kIFmbgLXEN4H7zMFDhgq7ZGznF1Ok/n8kojr6p8Yt4/yOed2aiFjqZ8GwxQ
Rtj9mpNfBPphIa1WP4ASKtXnE+IRRGXUice3Z2T1wvRtG6uOj/M/kZU/z7lg5t4NBviaVkQtb3iX
bCXZpmQTUctQZFbV9yTldE5Ib/d89OKxU/09uElnlzayXtm52PTc7oWPOqP+JF9By38Tn2MWH3ML
oSFDs7z2HdPkOkU70vQXx01LLDZbrPqr6eoJKMaPCjBG1O50+kmHGAzptnElRLd1JY+wZrXAhAxy
peg/PaR7Z2SRy1fNB6z5n5PLeHwFGdTR+bc2JYBb72nHq8S47AskhoEhOWnG4Mi0POl2K9cnNtcX
JeunrQQLhQkCoe2SlR8yUvITVHsOFMRQFMt3Oocyg1WyaRhdbmb+EZpswOQckx3muPR0VcycLpZA
k1pwUgRL/OItBRVtI8ctEwpP2w6IT70rnKHUpTrtE5/9zwIVINu0chM/MvPYEtelGkzKyX5v4WXA
9cYuqcjTXGaH38JtOPBaQRNs/V4Lts81gpkBHf3yMRkr8a+U4/fzeteLP/Yvm3Zl3+0Ei3dXHPOO
y4pOrnz1MQsrhm3kwrGAHby+pqWDCC0JfcDY4SZ7fR/9j+Eles5Eh+qdHdX5IEgCYsUFQzx/a/Rf
tT0JiWMABNj6RaqG1T/FFOQUhl+kJXeChggyTmIzVW3zBFajIlvkaWQ4q0p2ZaUvHTVvi0R0lBjU
86rh8NylF0grigbrLCVQTZ6P9q7oCzxWLDyaz6WFTtwydoSYtm39OVv7s3eq9Bi8Mr4x0h8pV4qj
HFygRopc/1KiF2OW6boUU5Gx2Rn1T+gr8OnF55V200mP8+UQwdxsB7AY0HLi2LZAtMmyQIJOIjWj
f1kTcQrj+/tCdkxK26/AGE0JWymnuHHxkW+GMnhMHZchZ00zewj6n6dIJivQWeWKYlB0BqCUEY22
xISK5KThv1JPlMvrDAsrXvkv/JnlZ5U48WLU/zY/m2+/7QVvK+vd4uBXkokFDpw14+4hBFODW020
kYpPJLkY0qb/wAQYsr77Uu+KZ30zOnZvyL8HqBtUJMmMpOYKTIPXu2nP4xZvPPZGKcojGBTvXgyu
eq6hVmJxR5sksxUbR6AXZ800Hr/LxBO6p03zBL8iAwRIEnv7YbqI9E5cBasTfjYm6Ne695WtxgC/
W7Q72k08uFihL0QC2sOOMabxBSUv+cXQyjPSLMH9VOzl6mvCTx/xEDaslmRrB13rV0HzijVuaPae
trlORIPdlWcVho3NBKVEqzBybH4mOnt+Ief5Z/Y4dth4Mk5gMhWT98qPXPd1jFKzR5yzvaC22T8w
1aWIjhymWZlMoU2qgf2H3g09v21RmG3VETPo88jAMzfOLJSAMaPTb4KWQwgAR5vlBLBWA185Sejw
1EO/xrZHuln2MJoVoei8yH7Mz5sy6eP+RGMzzDGjkBO+nHy7707xmRpzvUwgRMTS8PcaDLR0K4z7
VP0ZNd5gwS4M0eUMxQGSIDJVEKjgt+Er0aax1HJDr5N951EoCtTZ/Boj4hWW4Gm0hFyREsTrkVLW
3LmOVbljEHvO2RB6St1kBPpjp4faZG2V/5/E0ERtVD2HkcdLUasUL782+zuuh8fbfvGkNHWjoR7O
CYXGCVmhK78RhRnRcXHOyIftI66KrP6xQAwt/vC+ylOnYIBUko/Gzcbs6XJqpRJcIEroaQxrZdp2
0gyfu8C5yzbg7VEZ9PQc/G7lFilfGd71TSAqtzq7+UtqhRHeb4LB5aSDzojjrvjxjrDwtrRgK5qP
1lCNqYxF0jYhBN2WCGN+a7idb1VL7IretFDNZeZ3YiSN6o7050hNzO2sujxDxH5h5UGYkFv+qom5
P20dibyBRfCXb312BaO/PPylfNV8vNtGW2R+gipjLA1saPC8m9C8MXk0nbAbjEFhpeu/GVqQ+gJx
PcwZLMp873PtIy/eSm8K01uUTzx2Bu71zFS0uMFqet/gwbPfTY+U5oe8DoLP988X1MxwffhqzTEK
I/L1ppQRrSF/yvzpBnk0lyv5uOirpC8ZjUlSWpGU/XH6GFgJc4c8uwcHghEcE3Blp/FMabKgh2eB
4bJhhh6x3A8NCWUc2HrOYswP/NEm0r+leIZWfi3Eo0Gnndx+FI9szBWqMnCXyot5AmkLX3hk7bIT
y8n1ycs9esGQ8L/o91Duik9W+gyeMoTUgbNHmV8No0j6blGI34RVzwxbZGf959W5Ki+DA4yoJg+Y
EEbNnSXNPwUNqkNVIJ0B+V1LRccJ01C4nuRaHksALwNIlJrbmi4n00igf6PQ65BD86PFmRVMzCd/
1wR+8bf6rD4ibD5rfZPfxxzaCf1RSp7zbPEDAYQCbyptB1LirO+4dUC9C6vPg6RkSdDg+dGIoTQ7
gsDAZRIbRgen7qZWB9Avy7jsXVuMS4njMPmjSI0NzOU+257IbNsnD+XstIr4lnprmZdhQ0XkZsF5
g1pAUJr+myC66kP7FLr4ORRLDbS9MhLO7dH3kp0oENP9Ijeu3PpZhfBxVu7ZWZvsx4zBfchjqjXD
VvbMHjedvlqFSV7PyfZiBhtMByynFGNqP/tCEvfErtupKC+9u8N+PBJvSP4OuUjTzppt1P7NUSA+
JOQP55GBj9oCZjtAJ8KgDigLjGaXVMsq1I+DdpT8AVyF7ww2jeE+mH9yfQgM0ooL/s5ZEPk489Ow
8GPOd3E36e9/iNS/JT8dD68rCR2G30gL4wmmAo9X+BMcUtCeS38FogYhbsOGjsXDtvCUd1f4QgdB
zzCNv5udCUERmyu1zaAm69Et3fqXMHRtjmpBKM070X7dwwxYu1kRr6gZ6s9QMLofaVCxOcVRIvV7
oRoH6dF7CuGcOq5rejGGhDAc2MK2cWlmtMfYE8H2esypgmuYv0sP2l9YS86MZrIcM1ph1UrFC9gj
geHHcEkFL7QNR66foZEcvLnfeKGvdIollhM1oY4bG/q/QRNlmN9lfOF94EdaoA/REkSlK3DHvfJd
kL5o4UHzo2eeKALnOZO7gH6cqhfufmhIK1byXwbPbJnuYTbVzo33qw/RstCi/hslybyUfxZ8gh+T
eUzHrLnnXrKDw3qMgiXY34m9sgbHUgH1/rjIYKt4WcKutnvdy1Un8o7upseCslwlWEWoYDYT3lOr
TsVPJreiRBfBSoqwaNDbrrRxUNB4+9vraeSU9hNz683p85TKXysVRHwGG/PB+Mrjiyyiey5s6BGO
dicFehDhHgGEBntjSO+VJvkt9tYJRrJ+DPl+FIqBx/se6gEjEe2vP9X05LUU4vLK0HmuTf+5TGAW
zLLigvgeVnK/UXT8DpPaXp6vXlid4agKdy/joQL5e7HkC2cXqk8jDtsLwRVoiKqJR5F8KjSqPNAe
eIY6W5Tms3JNi1ButfzEKA9JXLfMs//LKmykcxzKNK/b0vgZvEtAG2WrlbEfpsusbwt923cnVBvg
2ldgD5WsIG1B2x/xT2fZMEZ0jG1/a0G84QL5CP/DaRwFVtu/eeOBlswWHQaXMSsmlFcv0UdP560u
1U1073NOOmfiDEbYBUu+JT46qhG3RmlqLViVEgvqI/Pa2zO2T+Tj55SmGCNzn7T6/9ue9av0D30r
jklhSV93KSgx4FWWdaO1l7T41Kwrzjz/sPSO/aR24OY2NcZ8rUJuIjebeZJa9CKmH4sVqvQBT/Ev
U9T4lMtG+jYb+oZnI9cOaqRTAnMhhVf/dyqH10KH8k6rpuRS9oPHBTqPWDo5EBaXEulgrNksJOAy
VZIRUn4Ko3dd1vVob4etCGCG27VR4x5Vgy+a3r6a9nQj7uW/exXuNCcp1jVU8JuEHIleZ27/ayMi
qrKm5MBOofn2WkXT1IjQN3w+BC1TzPNIsF0xx8AUQUlFKfDHnOuM/J5r+hDe8bOUYFKMX6y+FEar
grnxWU/9TIOPwgVetG9EYrmugMASU4hCLfLTi/OVwaIFxT1amQU1PltuH687VzNHSNlErQenB9Fa
EhSewphd5lhHFmqI+1MXZOq7423SS5MoMvkFRvjgbtWSMSihstddB3Whu+xpuFN1nVM7FNZmMDLM
OS0smuuFm9PlSpRmCModd19lqMiC+41d+CtmpgDz/c90YU0Q/aY+dVFtyC9JIwvxHPHD+IJnZHWd
ov5FnhGZtdCf8hlHzsq2/4ov7emo1kwRkfkQJR/Cy3EgYWD/rT/M2q9jI2y+jMX8WzPMg2rY5gwN
jBgbRsjpw/ADa7xKOFwKcILhizhLfPIQ2hDOOZr1aAmcTFwbzzHcbfEjKA2tpIsBsbBuUvR1JRMV
iA4S1DWFWX/65QlKKFyndobnKTi8nfaWE3aTS4dD3xrnp0G2L3b8ov6QnDzJHKCbWTeSVd6Tq76a
7ugpfCKqg5s6BmTbTOW1KH9FOlIQu05TCMeL8xo9+i6qWi2wqXN+4HicipBsZnLHbzw/GG+qez1k
PxXJcJ+shurjZZXXZfmyiBqOpXvRSOOpfcysJ+z7tVovSeFTSROo8kv63Hg5W8UA7y2jczP7jjah
1Emih+ZJlcnvvfZ9MucPlaZVo8sPnIHcKmtqdLeMTON+AujDz7W59Zur+XrYmNlT9e9rYI7R8qX1
JENXD/q/CnYXn77NLDvqq+1aF3xED4TMdH03f6Ig7AWKCFoh0+XU3GZG54M35xsafIoC7jXx5cHz
kAB++AY4+TbKty/lOg7RFn9ANRsKpimAhbaNIHOwBKBqDS/iiYUb8p6rsL7+Og1kJlqOG4jMlgDl
giD59RttXUEIjUSTu+z7d2wLGft6TwDSl2plJ8E0lO12aPr/T58cWcQlNFgxaBcplEnsfIMRWnng
5AZ+KRX6okxnFSPUi3jyhqJs4ojYbeVRQ2DJKBtUfd95N8RnvpTyhfD3sUIVoLbaW6JUYxndNZiV
mnDNeEegqQ4mFbQ3T5+1EhONHdroPYKS2/fbH0opkC0ECGBeHSVoJkV3DT13U6kNiesLnwnh2Fdx
YE9gi3InpYeWibPxxnKvOyCu4oe1H20vKzBMhgxGEu+Mhm4pTcTjXxYZ97qsdkYRdgrKHy93TXlE
nByJvmD914uS/6dLHmv0VtQdhCZamRduTwJypSROxbj6poqWc80rkG/vFWx0MvkwclRaAfBNbWob
6NY2pgDkNpQoasbVbYlOmZuxoXsOuKJbNKNrYkvf2IA4k/TjlQfgX1lxdN1NnqDOr0wSaEoVLlVg
94dWtkoL7A2iH7Q0QIz7Jy/qYpNYKaXujYxxo7waVzJlL/5ExYdu2rY45nQ6+MnC4W7uhJGUyMU1
VvD9SjWLlZIiTjkm2BxjtZ6zSZ9RxqM+ME7qz0H/zDYGqcbeP9feOzioYsd7BMqJWWjQu1YquY+M
ARkZgrM/qN2LQ4LWVJOjVYDej/YMWiL99s3xr/OWCjIUHAaJc8w6ITcp6EU5sCalBdrtPneQD3tE
lhi0Zmh/HsO48MyCtZqYMig3fyGIzSHXWeIZ1cGu2QShdLx6TeJMePX7DSBVkZWGHJqc0E7IEi/w
cERx2ditxzs+d2b8R1BIR4EBxbKPskdj7SdD7g6625en/WSxkIkl5DfZDcvC28H8rwS880j6Cybq
e0L0CQI8IzD7Kx/faUeh3h7Vl6174Yw0EE/Ct52cFIYHc0vax+s823RYZBUUkoyw7QwtDsyHK91D
sEFjV7fa4IzvV4IvCc5GygOHm9kOEAvQY4QbW9AnrBpquogiuMDeG5UHXIge+lY/4Pf/w14kzLoM
jVePV3Drmc1Kmi3yjPIqZHNhVN8aEzsN9edcplT43Sk+8WYtOYNXdSPvYPq5ZvF4d8POWXY0K6HI
Dt34sMPL2IcOu7kwSBAWnKDgwWuKGZdzaOMKbVr/P1sLz7p9Stojf4aKNoNrEexgaQoFm6J6rf9p
Qhcj9M9+buD89UiZXJ197l6DW/F7mJHehlGBgva79gdOanHdw5VnOdIFLbWtJQyI/jIJJyzFRb9/
nrb6labFSfh5wh+TU9MRG9z82Mglm5ILPELuK8uPfDXh7e0b8o9Yf2CmSBLEMrDst+NyNV4mnBlo
92USkkS49mISCcnnwvUePFf9wdvHzXV5YnvIxZQQETWn+FTFGDGlzNcZ+to2fFkyo+Zl8fD8E3QA
wdusInJ1jIHI0eXCKcSDqYob1GEoyqU5IPQfqL/aTfaszufDfRXVOQs4x1Rafo3aihPqYPELAvLX
QYtKOl8Ud5XurvOjsrZ/iV7NqMnkK/NHw3RKhhmeugF7RL7qG6b3ue9o/QYlRjHhzyxqIDzWZ7aV
wr32AP6KY58HlTwt9B6DDM7iGKFQqXrRqLU+j4Fm107vMAQXBtLOZTzqVc4ABXvlA6VPn+oH+Kkd
hXtgsHDzvAui69i4epRnvEghcH2wQR+C9+pUaUJaGsmG68BbzU/J8/NcvWcdanz3niU+Ew9ZR4kk
/CqGWjnY4CBf8WQmdjONWTYpX7rvav253ut95xNXocbdbGdJK1djlGY7493YbS7QZNLCnzB9kupa
LmfP9BSuO6tQa7BcZ/O8+HVVoayFjGpt+p89sd/3mQJUcfIHWgYgVcdysBxiC0DgNWR/1+M3tz+N
XHlyfLFu2+OLrEPVNR3jpGHHGt4zdakT2lchgzD43ETtyi8C4NUi5x2q+SDAnskJPUHBkIu+ow5v
A2ocVLSv1hmQ2AodNs3fVbvtBvDvMudhNDXd+GbZsRSjrLCZaf4+HsB6UO9Ycd8Yqff9eCwEWj8j
0LDru+mjUta2biXNbLeMJAOa+pu5P/Q672F0EqJJL6D5dAYjPrD0yzt3sx6eWFJfpJ89lbSNiyZK
69DmiyHzF/0ZOXcWCzOu7iBnrW1DjyyEXTu/Kc5YhCSS+qQYuxfP1KzWMJ67Hu0HDCFj5pe9RkH0
O5wvc8OcxmrRqpm3R/DagfFcYxPUUHFyGT/XtloZ1MaW379GZ9Cp8Tgv5Q7pH5/8EdId9jTTAUIf
dzWTJKaRBQdEoxaZbk2AeWXE8lpUVz7UCyMqWIEwK/B/MsV5Y3IcSUvZNe6GZku2lbGo2hmNqNCk
WUObxXnTaOcmBhxgLAm4qizbjjfxO/z4iCFDKD3VGtyqFXqUmH0cOenwZcovHgvzJXTXUiYF6d6G
uNWjnGJoxpj7xK1/CLlZhUxjTUoJQC1ui72K7ByBCEvF3Iw05p+lG4fmccXtkd0fQFcJ1kHoZD/5
bZ55RDaINcgw1hSvlcxCEG3IeBxfZBkF+H58CgenUZJWITPCEOsoL6YdU6rTxNNKgN9gdQyd4FmW
gJMhwy9/j1QoVI/zjKN4PJ7dV7GqCNZxCf0G5bdOYy+9gDRHVKWG4sgODYxXS4YSU4PBata/NdCK
7RpHtHozJ6nTV2ipzFMXxC7XKaVh6QsAQZsjgCCVe17vLtJz5skbtKuHNKc/rEtfUU/OLBJJWpZV
3+hYVLqxNCQc4YGthgXd/0sVa5e5rD7z2NpG0T0g7IgqznkP9jT91DTnrlB8tZVeg4dKVAF8Jtqd
ObYUlhuzxlxBtb7jnwhA/VrZ98Keg1p0/zePURkcCxFE913ZqBMn7cUe2CPiOGWVIPlFQp1K36rW
Jw+wUUcy9/8MBU37DYJyBtdpelNrRIDcBI4vt588oWSzGPhHqFSmABqf2YNn8EOS7xHK8YeFSKbR
DddL79KPmAPOuC9sHID5sP4i+jnhrZVv30vx5+8sM3MzeEPyvsyzAVaGubpJY0v1z/haaoXWpPwI
Sa1uAT+FEpULA3rosFrJATcZvzT6k1Krdc0kqjOwnqGqSP66+I1PfG1oQ0/BTtSZGd4/YP5JfE1t
JkoJ+/Lp4XuRAukduv865NfbGsGfzf/k7ahjSikVe8qWX938wD6g/62Ha5I5i6C9oqBAa0L04F2S
9BsTdUBQOff/9bEhhLIj2s9MH6xtDYa40NOXOhfT/V6U+jzO0llqOY2wEMakoFKJV/P1W8zwWcvN
9+4mhsp78UTIrpr0cw+xw7S8THW/sWV6NLSNSV9YHn8KeWEsRP6bzuqmxCUvXPyzsrZOuyQTyYgR
JWXBD4lb1QoEKvti5pdkPxS2EpRfuPs5YoXXxsrDcfLB0YdDg9lKl3/tmb9LJZVZ8PqHpTBYy1+M
l6Wbg5dpyPgA/Bv5cXBNNA2SjZ93w+HJ/cx3nX9vtegj1rS2Rl4sR6ty6VE6L8O6H2rLug4XWaPP
02LyoTGO1spomH9+BKMMwRoR1aquHLLCW5temQ59e3xTzryKfnBo6jW4RpvuPyRutZYVqe5WEON9
m6TbbFQSOTzu2vNufg3pvOn/0+wcgXcwKK3T5vHMIrbt6lqSqpIz0CepwPnXLZFGOII1HTN+XWXA
P5glbVWMZ2PQ/TD34/Ky9EIhlJJRoy0j26KyAIIoDdY67UmkKyGQTbIh+8tlrYRgqAVLY4+4GEiQ
TYYEcYjBNqXSeFJ2mzSCceCGwlPDVhBbvfli7K6kUO5En4pR2rPhAMpolPnXoR1yRnzme8qGymy2
HaO+tmS8n4VGzzTzQWTVeICVGkPAJwfo4QGNC3URkXUnHIGDPeSZyJTFx55VM+RjKhFMmP29wKPf
/dSFF18uo/58Bb2VJH9Z33ly6MDsv7ob3bVdQCdJxwwRuF59xcjevMVPfoiF6kvtUWjkZEmKCCRL
DQlrp1ppScSRZhWhmeAn0C3bJEmWdLVMwOgxV7mr7WXlya9Cv8oPoCbh7yu/uRvDUGnaktXzJG+M
XidHoPzphNtMPCLSPU4qb5nEtqKPk940LC4BaTXZYjv/McxDkBNrlHonKv0MOr89KXD6WLTvPqPf
IifuyjpiyvDQ8GDujNPa55rimDWoqn97gc4ltdbM0zb/I2IJXyyHwKOTlatNlwPbfU/0hupyS0jR
bPhFuXca4c1eJCMbSLA4nfdKySKirnNUqfx1Gv3xaDO3g+5PLtBoK1A+rHahaOolBlFs363FZwXV
LvyUL+SohdpRzXBkL5dFKGOH908zSKv6BiyxScSrhCm4d5fqYAHDdgaZkH2zLmi2dPMnOU+4tt7a
fNJJ73bOknuunZ0L0lvFQPgI3g0cMDOUMUb1kYdcY/Yrot9cAapsh7JFfiqwP6FYy3MgTI49NeCP
6K9J2EfFIvVH46QeD+u/t33J+F5msK9TWaeZRwsPLZO6wo9osONRqmJggJkgoxbr6NHlm9qWiFan
ngTuOV9oWaK7Eli+evQ5PTpCzAioLdFTOju1SehvCVZxI+1PPbJzhk29h5Z2vHi09G8xYyoYNJf1
PG92e2uixCKsL35pAAtfryMzV/p5NRGQUwzFzB9AD0HUvTytq5wBaAXUnI0ohHasVPaTEZnYGdfH
FIS0gsVY2fHGeEAXwhLJmRCzaaUefN2o096YSWMvwkoR1wr4gZZNr86QCV9Z3miTqNQBAxRUdSo9
ToM2ff5JII0Ll5FYw6DG2XQRaZ/j2dgec9Bckh3imY7c0SLR9SGBOEGs+3EHtdwFFAeJ7FmM5jWk
fyHq6C508UGJaAJ2NfpshDlDYYPMHFLu9rZtmFcTYbilk4Vc8TwSzp4hlF1dwttYl/ewtH+TUpYK
jamOj2ru9+JsdSgfFq+0ZNAByfgm3zgqa5Pb6kmzs+pGVphsA8hpldknn46EdRsZaUbY1CoapyoE
Qtq8S7zeKhmD81heXGPKB2XkFxr6nABLT814/cnbLK2DTglfZwMtGWoyDfFacG4nfGxpVbVdu2CF
Rz6vY3fBffDypRiEJwRu1ST73QLzaW6uC2hYi0QG25CMHBzs0DCYGwx+RAgIgXM3JA9OEH2DUyFv
u22G9XzjWYe/PapHRdgbvhIF5NZB3uVtsR+HH/IrjR4YP53oz9wJKSk066QL2WBcB2xudbqd9UlP
N3M2sucnE5Baumu7qNPmzMpvsMpZ9ia9H89/gwGIBtV+Pql31uh76KRXxQFKE0gfMRRR/9QFEzDf
6WHKkgDThAxpwEGLG3bkMZX/Ui0D/m3sbJpWLv+tjfWUvcmUp/l5sq1eHkWmdWDRz+YL359wyx4Z
b2zlGpVujPeOhEQOyZGwrdfg/dINi5i/oQGGKURTpufECPCaFQr2hUmsR9pTK4jGPNqsJpd5TcWa
a7ITpJZbz6ATQhJPWt3x4QjMc/AmzLdJhFDzxa/PZH7IDYccbkPcosFZlLuaSwn2mkMTwiFLAphO
ZoPpO2e3RU4+qtxY6GJBOBSk+9BPc07v9f3wk/IqwP5PDuG02+RKxEhmEO/NgBA41qpTUpT2szLp
7qQ+nifcI4NV4NdVZKyEHkwksAu2G2/SdfoQq5dW06Xj7OZkhChQYN+4okfCm2yKE9YteaxOAQUu
aDn/ygsKMu4ne3d5zfR9yAfS5aJDez7xpBSMMD2yyoOx2ZEu7D3/GgtfLmmtfA1rRH47pCqzUaSM
jWmH7WxcivD3/NWlyU4D+geR1FNaWfOCpMTdqCoP1x979VRPs0hWcfrF7yFNeprXa1x14kOshLDU
I27VfCVjwbq/hbmEMntuAabxWpeFhgOmnUL2kyrmM9GPr6iwrmlO7liZcEzJ3O/eHipMXWVYV7iU
DkSOR/CQtFcjF7tCPphnB4CnvB17hzKNqM3fv7mPqC/+5TCauENIDiACgYlEfg3D4FG9dMb2nYP8
avL8AH1W6CUKt6fQL7bAZIw16xgEEECfrK0IJlvPR2C/qv1VKaPVcAP/dq42Vut2gp/G0QC62PAs
QdNU6Uwta/RyX/ZG77hFO14ECC2W3iYafdAzWHXs6rJSTfnEwcTlPNsZkp4ZkC3mm5f80yRUssqd
BHhokjL6RbRXvHypYuiiaYz7xkYF4bab7INXiy4wCzL0c/iPRIQd/+BxNEzQqmieYLPkbmC4j+rJ
Cxm5fQaUqPxex8S4yaXMpmPYY73Cv4e/P68aLJReREOyLkx4tcfNUE2Cmca82mJj0UwoTUGYRShL
N3RWpPSJDshJsPNFWZJcZIpKQxEr/CAS9nro5sP309sAGqwzRYJoIZavVYNE59UJcLvH39vtRbFb
krHgbPCt3tBve/+vBsR6NM8e8Dx7T3Kok7GtNa+ZReSw0w/s/Wbg+YTjmSsFeM9LKLRTctVW7Inj
FKyuoNG1IzDXJgHIoZqesDivotsaphCu0fUvKi08XOB3ri/ybAH1kRk5rck/SSHmBtB8/sIvgG6Y
w8Dlpb8fazzNJBhL1+YwbB93CItDVRYmAvXFwihnVlkqCkmzjyMvxYjpZqrvq/O2qlawK+r6yUO5
R23MbJWNzd2QndwkVfrBhVg8YxzsVJpCRAvns8iN8DVa/JDKl9Xn2rawsob16QSt0KRKdw73WylA
7CVZSp14AND0m3scgj5/aaZkodspLswlq9VE7w1gf/daEb8vUTMQTJbSEtrwCcvc6SxXDbc9g5di
9cltKYPvaWfH5Od314eXPrvWqbB3t1lZkYLbXH3PmAcy6FIelqQ+kYK5CfehVHkMZ8uZKpuAa82F
aLPY0WuPQNnH42FF1NbaAFL/vOBH8Z4a7A9O+SDRr81d0qlVR09CpiF/0L18GOvFz5C2ZfFoghpy
qGrRvsnbfbYVO9Z9OFMoRLqfZlfzgWwcv3ivYfQM546KpuMWchnz3ehmda13pdGTN9eLBu+olt+k
zC7sUYpGFfW0HaJmYUe/eEVM1R942uRgBnHA05GL/NWz0BVmrWowldb+DPVZVTJxDjXIpp2pywqP
t+h8ouZpBjYOmlQjpCPG0hVxCEVsI8Ac2g+s8GoIZUM2/5m8MnpX25y6x8L3VKWVcsw/SAW0bR9u
TVoUsiobNrAGBrs4DFVaBmkeP0lArD/9gzJIU52TYJ3i3CLjyGvlagODJkMgHGzUwW19nJgLXmcr
iMXuM/On1NvMB1q99sIIbzUSfpxrtdSlFiZhHWWGTsVpVOHFNflyBGjJA05HJct/eDcNJzSCQOlx
eQn17CuQMkzjmQWjePgJgLGS6XrBCFqHGlaKSm2Gm6pxRA8w8D4FhtjvUnNiXiCIsExyJnBmYapq
f+rP+25VW6oX1DcGAoGjetsLXAx4aq2GdkuVNlYzz4TRQ6Q+gYBTXnh8DFT16fGEhja67ihV9xP7
yTHBp94jlMQzqF5bRrCrAkttcrqtPEDHImb/0M3OF5v1jZnGu7PhfM3UEH25Tk59tJYqZJtoe8VI
yVQhCRlj38vkXJ1Fwqyz3zPpFJfpXbVZiYs6ry7j3NHzzye3IPWbPSkggCL9QMiijAEDhLtWKTLX
u5J/JWBnRyJ5/ldbdJxUR42UfmDAYRTyu5mRDmUTwv84ofw1JFZPn4Sv7eAzRGBXTcLSN8yXq6wf
Xs7sym4JcH1oZCfwzFxmC9gHK6ZclAJACSe9Ed4WJwrV5v9AeDe3xMrqaKdXgeQjLk3/1etKERvz
N5oucCJhNxPK6d69RqzQ+XZqml7NVy0JSteBESG4AbJ2ZOyQa4OUJuwtQxfvb6/PBgjXqr9zBFDf
pzT4zMDg1DYOy2FOJkIgnmO04gYvkfePbXrO/TbU+AR38a7aPqAEIWens8R/JlRVyJWT2SGULjPr
kNvyuN5M5mxCrloHpNOW5ubtUpCLhugEwO5mf8pWd+OH/Wfa/U+4fcSUNeYCcVhHXHrUuP+tkKFo
GMyseAOC3se9UxJ/NuzLV+yhob8z2wZfW2iSeIa4MiV462slnVWmQd/NJRec2kHH90qtB1cLFmIb
MW3rVAlPCukcwnqE4A4G4tkskletK+SubLzgEiW1svRIFYZoSc/KKrNAlbBfThtEz+snAW4qwEUs
59Kvby0aNdvOwj/axvC3c6KJ46nNLod78WI1la1ZUkhlBpFEWYDk3QSslykA27Yuzj41RBO1Yrpo
m0Iv6Htipg+NsNypPjrc5VSF1q5xSkY4Sq1J019dlaZpLjguGtBebkaKVzUXCf1PymHWRndpaJ/S
qVACI8qQT7ZfaCW00XAqXd+2i32yvZqMfxvE0N5JJETg53uBNYPicfG+Aky6Q7FOkSlOV/qClGIr
7oYPAoszcwtOqs2QcSt9ZPk4knAVOSw7VngxvGgADZeeCJS37WHjvgwBQrWCzEimsT6EjsSTY5ip
cP479LL0jnJmcFZv+5dxi3QJxQqCSHRzyPBI+hPwSJb4ntzx2/G62O4N7ZRFE4C6PNF2TETe4z1x
oDBMeso9aZragtoQ7o0WXG+Y+KGQPBnExspuiV7OqlR5YqS5kHP9791EBKKLBTpqn7xxFqbCY6rU
BxjA8JTRU0uCslys5gjB6QQoNA0Ot69RKGFXX6ocrE5G4zglj2LL0zypZXVIV+4+ixMhDiCTWsao
6OWZ757KRBV71PcbqgEpfAWHbmomPBAY2POOB80oyi1vumUZiDsUD96z/BOfxySXZX7ue/TQEo4o
+JQop3WBwrAgla/fA1HOTAxAITtecA8BEySVSzyuSoqW/pL87UDTsne9FuUWcCgS9+7eEWTzlkkw
tPJQGdCElMgcm7h/n0kqDV63B0pVNa22cxrkUJ5f/vf31NMCFDpH2yslh/Qvs2FNpzeFd3lKeRTF
vRD8shNk0ZaSEgTmpoetesPjvhzx1YPyxxmH66XOp0bZhBBGlROjyaIrhb9APNuCPy53YTNFq7b/
LAl+1l8eTEz4XSOpImdQpPcYaXaMhTEr531Q58iT7+rYPc0c9xTwWx0QtNw0juEI9ZEv9o1oLqVa
bar0UoeWBDqawMPf9eR4TerSRF/v3iWdEL8oWLpZ+rLja22ZvtTopO5eS6Ejzf7qdcInc7enfgjU
2SGDBfNTBDaAB+de1LI1vOenmh7GPxrcMHCejRb8Y5PeFxHQbcfj1adRr9KKUN7MgD9MjVo4Dm5Q
bm7XXreD7zXai7Z9kG8HEhBGxg2vIZfRnrnMfEt6PuEXNSEIwVOBAmYsY3GpuRkfLBZgA+91UL1P
XlpF/ic/oC6FtcH4Ywm1W6doZxX3TxkpAm45Uw4F4MNpDv3JXqmq/zr9+xmzWCZVDSUVam0J0PLH
H422GM/iX48cXJSpBTrqL71D8qZXz941udhLeCo/JtDAvdto4GZv9im5Lujrco6Nido/PHE+S4Ii
62pJL9OLC2wJj2FZ9sBJQZ6JhjTl63Tth4WRWa/SvV3Giad/VF9nUSDPtZpT2C8vF522c8Ojotke
zEyfcV/CGoJcJhJsAwBbWeP7bRRMcqTDJ6zQlKrQWtxsCGwV/yMZjTDxmDrAplO9v0SWyan17w/0
la/JTv7eYThkC1QaU+tLr6+AQXmKgKCOuDB/uRlcqYdN3pknQufaSGvisPsMQNNaNLJ/PIMiVRKr
6VGMEMVWKgqNLVpQ8bCLtBzpwksyWYInhVHTxc3GyVVIQ4MZZuUoi54B4T42DOohX1rAbN7K3vgB
aWkT7wWJu6vd7miue3+wXIjKpe1Zo8x5m2OsMhvYTSYHwCj1VRrOhyhCyiPVysra2vxC5VNNNASg
Nj5hwboCEIMytzw7Grpo+Rhw6jwPZ/Q0h6oFEClzcftDV59K2NhgNXLAUTi+bv5GWoK8NPYjvadv
5gtPmdjB8zB54FcZcuUNykfaGwaPYBoUbZGLnJ6EYr1vdjSXkE+HcRC3Mj3aQOuM7bxRmMsVUErV
MhQ8jL6qG1IklsZqXQoQje73IhisREg0JflLXuJqcFx59akYuJAc2LdRZenbgkHVt/NyxH+h/ZlS
woWW32uF4cSyycBiYXRh6qXTxKWYFpqJcgQbQz2vwqvbfP13auMDZDn3ZWrFFfM0Z14iIgg92uro
sI6+z3WMgbGe7+zNOugQWldDfJary+OT0hkn9TuVBVL3ziH0H4R9D6gXRKklHEJLNEj2d7maY44X
3n9a5dsdEU4UAzq4AQZyocNqc97wHNh8tW5KAbfhmWNRTk9EDYRBSfRQxbQvqzzRXjLwzMieisox
WOU1h2lWkkgUcdbBttXEXUIGlWDFmUVmhAb5j40SMit2YwoIJAMhTiX+jfgcXwtJr7YoN81bu7Zp
VJADrjLxWokLLFSyyJ8nb1u+n1r+8CR/qcvXmZ1TIwZ+mVIs6zlsD+gOZAaUgrxw4z/s2hzS6yft
/FfN0ghIiS5kF674++GOvd+uxevsTmPV7Fv5EouazDFwEhql3zZl+PN7hQhdSq3DEzOOGwWvPRaR
Er4ktktIwZiJoypJ0q6PM9S8Z2n1yXTv1DGWbr0m2dRf0v9bsLvBk4Utj82sjM1GbqkYhSbORm2u
CVn7gHcISHtthGt04XJ01U+Q+EkV2cvg19F6GUjjGV+voV9m+REA5gmOba2iI1Y6aZEN59JRx3Xm
uKcs3BbIlbMZlNqoFpQO2NXYLVo0Z2b6aUTiWOcOnLNHbs++rVEyQr6wqudrNSuUGy3BJYPN7FRe
tRh7njOhI7oBzKp7+EiFxIrjs5uV+76Guku2/4/rmc8kb2SE4ggEuOi09Hiq3kKKRT6njfMCU1mL
o7ICHqfKoR4d+bpZeynGlEp4sDeG+DUt7cnK4LHvW7GiexwFOivBObTM/xVBlqcZIDaE2bIi7bdG
WoPc90oicdbROpV8OiEtaynmlh+5i4zro1u17kdoVIf3piK/qjiy04syGIFoLQvmSAO/1dUusr0h
t24CxMUeHg2LvScO8wGYdrolESlW9VW84FEPpKOq5ORvanxS2egHRfGeAdQLApzhKKrCIkCeuEC6
KtCO9euvZFu2EPm24kYq7xWjWZdPwBSItdE5HdGlN1JGQlqtxlvCFe5i5zJGgxlboAeAA1iYBeEo
NRzHWIXfbes5lZicoAQEv/NxVSP3H3uFZImvEcztHQzkIlE65MSdv0n6YP3CIIW0l5Omo5Y/RR+C
n58kvymQ+YmBLXBVVO4gT5LCoQsiSk4LgWKXKZhlevU/idUmTiFSdhzA0/IvF1xkoEVo2ccr6h0Z
BmGkCh+f2OtW5thHzPKO59mRwUYBO1ygn5aQ1hBA6Wnsht1YDDZenJoR8lXc/fO9/ahWR0tP8PSQ
Gh83sCmUnQ6y1fe9XD787YPu8tKez9epIMXS9eSvIDxTE/RMaoKL6BkfzKbHiH0WidYSb3EK2fKw
pGr4mEUN8YYi+woAesyQnxvNCFGmVL/j5bVd8ut2+AjNXPhoosMzWeX70BObOZi1AhCIQX707eKf
yDVfpbytetFdk4OMt0DKWYFItQfca+eLSXgC1OAdMsxgwU1Vq7uJgFR/eTo/07A0EKlksrJscrg1
8AqiGggKoYMgKJ0I/A0Q5SsR2vXhRhkY/7FtkLJ6KoQzDUxTVKU9yhsawd/TUm+jG+XzfAhRqbxv
jnErHemfOPcDufFYNBTVpWtXfceJxIiLqaoaDoxmhoeiJ/iUaia+inRc8jRmsJoVELUj0HuHtAQo
dSa4deQsMGTbRFY++miHgzh4DJVLT9poMHYXaL9kkBXkPXYsQ/BPLCDP3MboNAouL7rT1UrnIWOv
eMzUFFsuXuf4jcn3EOzQfr+bPnoFNgCrFQLYhH0speOFF1CLiMmc5HSpj2jLUYvUfr1iUdIww0tb
Kxi0s5B2mwiJRm3nxyKoEccL7n9D4H//XykkklwH1xVjYow0jwQ2RiQhEG432BBONY7SaZhKAO45
HRwRdBDisZpdptRc51w9pJWZbUPODmSSxT2zLC7Vkxiq54Gn+ec4wA/GOcnbBaVTtsqFGa5Q5mEz
LaayASZ9kVDtGIAksPighC4+qSlAkg3wPOWsji9xbLvEP5eUM/DfyIbe6ORTuynGyNycUdcot2Vx
cJgmbi+DeFIMVLzz3bU/Q6PrcVngItrshK/Y/mZaguwAczAmIOPqrjIrmnI7pt59+87pA8h31+9q
zjCDybpYYytUB/mhnBpMDhvjFklcdhtQBfAH7ThvBb+58dPwR3Y8c01MpsInJOopBaOjXH0E4Xr+
7wreJjuln+Zgam7eYdJi3bSvdS4/EAOprJ5cv8ciF6aRr5m3jwYQXyp3+lbgWI9tRa1ojMMrXW0t
ABI031TyAZjisZgtL5BuwKwnfLdKnhxJBrkDY9O/z3B0+/winIQRDPG7CFPCKu5R1KfGEXOrF4Ol
YoYipzcAohrX9KDxRABhS2A2aH8/F7fSqs4CnzzWBWp9+zUUnbwrfGjzM047hXS5SmsqhO7rnKpk
J/ra8m9cx94Ur1eaoABhkzSu1IIoikdMvPLdBnmhn98cJdvhi73xKyJrJmraCkfVSsjBzTfrxlGs
+L5eqiIybsDjN5zoYJw1cc8j6TYoAycVPmMAvF50K7SWSn/aBndIXpQFTkjbFgcykaahx36cVd90
KQ4zIxfmaUuMctA5rsgSFOrkoovu7w8iYr7uG/zFPQVDxzwSRBwNQGOoE8mvw3Jyb7KD9OnqmvB8
FtH0dIPrltzvVjidgZbvIfKCdkZt5sHPRagJmvSSbr1Qz0eOilFUPYeROTKoLq5X45+qZTgHwpJ2
4o+kfpx99RGbcNIMHit7q+u4eMD4vpGbVLjMV2iEbTwjnqYQBGgEOD4EKAwqDxWWkBau+/CCW7il
SHzyvLJNXYXbGW2k4+XcgMsZ0lmgcTXImfwoiIT8e4eJtWocHGp3+HvIPkjP8rgLDJxErlapf42V
6aKQOdlmPRJg1ndk1GC4k6I+1nroKQmfbNh72heJDQ0x/XmDkASYYlyUjmLtIFw1C+/kgXDWdKcH
O+RtiSodHlYh86wZG2UEboOmVjGDKfBZyLYvWHpmuafhUb4LABXiurc9FyVIR5gnug+3PS2Jv/ga
2ABuNwaYf2eu8G7gW2+J/0y4S8VaZfxQ6IlnR+0lxhDxjsXqz7MeCl4H91sNMz0LPiCkNGFDlENJ
8po6s2PhN5NuxJPTHNbJYhf7bRJlWxyJh/rWm5rUIQfbUCMWnrv5cKhk0imc4IP2Mij431Uvl/KE
X2pnVCFxcCHDSNDCxaWCphiIC5MHY65ISG8fCxfJqzzk/bBK3r/QOnir8icnmLRE+gjhvyt9EfHO
DWJ0kKtljZAKuPFsbTYHlEx5JGLrTe1L+MWd2GUL9NzqLwtI0T3Mab0Xf9HNGqif0p2m30a6reMd
aSiTnUopUH+gPvqtcrFQWlFyRiPYEIqidQ82dTHUjiTjALnvZdiY9ytn95Otby+WneodvcdkAEEB
p48SWGFaYm1dmCjILYqucPVovXQLe3JEheLSVhhlOvNZYQJMagopnPOBNJHr+7ZdgyyYHPmxR6ng
3BI0SIoHmFVv17Ib1LzAIBIDRoCKUYdVLKRrd2zL7UHbpv/SocwHtZ1P6izHbmbUSXv8OL5iENm3
zYkFLAvCTCuPl3E5wDOI9CRUVvUlFzjcqS9hWqXpdJOi5xWg0Rj9ne0xHOwbOCv69kaJAWVDFlwW
BC/KscXKq+J6k4EHw/uBE8I8oxh38byggJ+FW5/Gh9Wf/Ifdbu+wyWpTOpIhba97WPdnTPl+fjl/
vI6voerhIJ29zrEnsbJS/lBzQLp5KQrfbbJu6rj78C6dht3J+XxKYRMIQIPplPScAarTzo0Eqfmq
tLNp2g29CuL4+D2vxUT4Gnn6vPJRoLAaDWvMzSsyxdJRuCLa5fHpE+z2+fMMYEBld5qkDKExDnXn
vIdN29TStOyum8q4gbo2TcPPvEXSW3UeUQcF/ajhpESQYCkDB3YdTyacCNJOOXh4KlIVEApl9yBg
8cISLn4bOVYQIBpV7ReSg5ADZRWJ+gRfJLcCM/FPdRhFvyuCoIBxxHUiKgbXB+EbzvrWYA/GAwON
plS5xWU8LjaxUUiR3Xia1WlI7YAaO348aTHGNJSH9jlAxAxE7VfPj5ULxT04ySJdrw4hMq4ZTNHI
/8s0a7rk0mxM6t1oX+MRj3Ep23nGp2gqGAqt4E7TzIuyw2PZE3Hbx6Xj1cu98kQK17ewHxR1nB1e
l2CXNtGRIpgGfl7j8hMjdF3HwuK/EvSC/oABH554+iY/Zg5FNVeY2w6Dc8cFMx/TQdNwqBSxu0IF
+3dn4lnwJQagzFcX9z4X9JzYzT0z6dDjfMKy4+w+n4dYOm2Ag7ISCI0Ez7LbL1AMK9UkEtYR+DkW
VuUXLpZzeOAZoN/v/TxraXwhqvqW7392FwGZrr5qy2UjVU0UApFlNjszLZmpJpem4JZ9MtOfwdu1
MGahIAMSE8AJE8XcqWdG2A1WYsKhv0uEaIlcaPq0j1MQs5XDOgxMcuyA9QWzZgBDO6jCFxWGubIX
ulzXT1Ky9NR2L2kbTjd/PNp2UVT0/tsjrrdOaU5bJ5LQ1TO61MqTn+/pa50o3w/NJOGbKr0zL6Ji
j51yiGhogqFb3W0+iqII3aDT0Pq86+O01W3xLYJMfUOSzFlPdl9z2Upimd2LfJMlkNUGdl7fHhCB
sCfRKdLXMfh/J6p9VcQ90GR81h8BD4jcxFMnD40x64ROszfc+NKhOHHmAAeZqm1I7fiQ1oHFX2Un
wVjniaQo7LYGt3T1hNycRCPsk9llUaI/iTgRFXtFngtSiefYufi24p5qSvtMKRmk2vV2NcBwefZ2
90AOygnhGEOeu87ysXym6QoiV+F42wtS5rMUHpvbAqMnTjlyJR6dy9YFuH90DokojYIxmH5PrgPd
88J3NetGMx90IhmwWCcQC1MChe1vpzp8Gfqo5lUTKgICvYREC49I0qwA8kMfoKCFXgg7GnlAu18T
ZrV5xm89zkOCiRbw5UEJeeNcNLiXHZR0b7Zv0jKyR/IgCPIBfc1nXfTB1PZe4hqhxAjlBm6UOnCf
vqJsASSQ7vP5Fad04uvZj8EF06piBCJsQSD5F7dyzi6n8sOrdZ/aOrDyTULwjjjTgfl1MCi9enP6
9umqfIE6jLxs3SIOckF+n0+cyeUfW2GHvkDz/P973ZH+4zeZgiu8671YAEZJHexh0Ezhmly/BKaD
GWPKv36UEgg4wmpSxA7snDJaiBay11IZHjUSXnqqCnkNMPASBTkIpS0vh13hIIPtG46CBb43Ewex
ptSospUWj6rlGGuZh27J2Oi8l8n1zDXXqnmBOfrFxZp8A7/DP1JjSt7U2vx50F8FPoQ3t9FbFDjH
rdI69tAiAwcyKA0QQOCu1lWxU0LA9aBWuRwTYOucBdNrBKi8/g7uI5o99dSK3AtoezYHb3lFCJvU
kmwLIC58N++oPHDAi3NQ5277iv6OtyMoLGeYzJ81fK7VnVabBVXYk2EqvCl6SjKMXKtseDFB2VEP
DHa+0u1VApg1IC7Yc9wQ3qquj45dkw+I8v31y0U1lp+xp9wOayUHdN0YkeIg6z0s2/joOSXZyKVw
hXYbO3vcO7VQ7Mn/rksS3uh3Qu/loBcfdd3q2H+8aG7po78CrIwEqqmWaJJpO4EhvVqz8gXKSlLj
bRqtVScw8FhqKeK4pUP4ZJOL+NoFG8RGdyUzA3JV398EjeRPxFuzp5k1DtRGEJVPczTm7yIAsl3I
OcE/aEFA1CtzjTg6txu795p5CFFDdtX/pD5JaWgEOU4YYhcRddh6zLs3Eo2EMmCcDVr0fj9Y0twS
doo7jCTFT3Mr/NyLcS8cUcY0L6XUXFom50WQ0OWEB7smxDuWqlrxkShiY3QGwQx5X72l8AalDV5T
9UCbM+lJLsWQz+v9VsWX7XP11+f8++Q2+M4hXyjFzT5cF6V6G4JOlZ9RhIOCYkGFCzJMO90e4DE8
Tm7nSZHMTwjy6KWnJt8qzNYCrTOrrCc7hNBAhyXwbl3pj2CqnJ1o83Pcpq+vvCtfuHqPeHt4AVQb
FpnEyUVR4Cw1qlWPW1c1rAw5K81P4DxuJP3GrSfrL/lEtfToCsyOIxv4sWEP3Sv0ccxBmitP7wj2
qd42aj0Jo5PQwxK829xiahYLjLkNqp2WJoN+fAYuI8Nxv6s4WgQoTxfP9IOQYAxC/H6vMj7h8meZ
rJZa5Zkgl9yEF8vDY2nCdwaFhCoTny2OsAPoC/DrO/mBZ8Tqsg/oyqDgN0xymyYxOBBQTTQTyvdP
drEZH3/TPtIUVsl0Slhz6IXQFuxzfp1tJ634JTyGAUZ9wODJtOT+EURL1LmymGsnRlE31IdlSnu7
/7k2lJqNuXTsjeaCs0hDBk7NAl9EzXvPnBC24Nq879DHSZMi3wzasCoERcszmBi+mMG/A0TuCBuU
ZmAgB0DezQjQvKQLOgpQ2JjBazvpUPPbYnIbo5yPDN7k0DA2T0sZP6wXDl8j2IcXgqhZob+NbJOK
zE93aG8EuuloemHhSTTt1gAJVpbDjsJJWFbULo3mUm7Rz7m+sY7uK1cIhytfXEHD76yRSzcVTxkI
7FzMivmHdmlHylkDlkzyGRch8PbtIy90CLEJwpdCYTJVvduHmIZROvYhwq+9YYXRrNlI2Gc7//VZ
2iqCG5QM8z9wNaNYs7VkrMxMuB+HeL7RrQ49mnzOzd2okaRTIhWxErRqu3fqXbabtOf2u1HQT9QF
SFopobnCtHEGWEnIBo/WxMPCAmIAXmx3qbf6bmLFUFN3ypmkvYbRB2tMM2LJsNNH5nDy1VwjGvl4
iClmvSUYZliHsLxCYs71u6NbfM5vOE5tlZE/sWtjczsavKkvMn6oT8CjKD+0igVRVgOXo9kwtD1V
BUTLAxXDCGfYyedXAbFjpyM4WCkfrVjB8RM7RiU1RN0hM/6c9RqKniGW9Mrvou+mbpkYzqMKqXY0
8IsoIV6JzAJ3GHPsUfrEno5HQ1j7jy2HQH5+pXKkO71xoEEtHnrLCk8AkskiDA1BQIH3njTdK+fZ
wDI+a2ZM9JD7ldWhobBFPV7EATqQD9UbOww8ecGLZxX6d7+ssXI2g71o3K7ycnHwJa9gjub3TlO8
6JvDSd7SuSuTNOPSR6xPQFKunOsOp5Uil+hJDxuYQk6TuppIZVCABwkl6cjhLpXQez7nH7p66vAA
atVK8lGbkLm3uBOkSEHflBuz9F52+O58j9RKX1PUWOLTQ1g4NXoBg/DADPho/ELZipZo0eE0hX8c
7rN3DZ0LJPns+2+Fw68vV2curPXWmTy9crqE6VXJqBNZ/TVQwa1/j0PCK4XOyIe3ycNFummHkJtJ
h2O5M3cDbKhNraWnY7BZ4pNpkp+rqTEdtR7SrXukxJAC4ChPXkRPst+NLnq8DR3NIaVNFNxBo3cU
D2NcSWAXU93OmuKakQx+dEYpg8Q4Jkb73kU6yl6JffXhIBZomz5cxg45VIZoWae8xv9NmeN2ut5a
chIeE97uR4z1Kgxq8Ao86U9KRYOiSYSpfwu41Rij5H4h/Wbtv0G4jWw/KQt+dE+15UaimhMZAuzO
iZ31gwOTw2RI0D4PFlDzFfUMSMwax0P2xfLcLk+8C272mPNDPZ3ZbI2u6M8Tz5+dxEbujUSyWjsa
FpXSKy9MJetvtfiQyBZPtCkFOFb0PWBcigZSpTlKK9p4+VwtJ4cY49pNxWA8cgbgwedZJUvX65c6
99dkrojpsDETzdvEQXJqr3A5tCn3jrhsNVksXzbFooKnuQIZAScZgNHKSgcwqBwAtMx2UGdoncVz
m214J2sRzDqfj484Kco/nuEQx3g21IfpGepol3Zqn5Nx/8AZVDZvE5Zm2/JIQjUOX/5q1XeD0Ibv
Z+d/dj7zVpKVDryKW496k+aoE/H9Zx3ms0SNenEz/Hrfct9xTk331jlpkQ/pLSaay1qciS690Zs8
Hts9mEOMbLwTiRM4FWb7SvP9LEgheUzG44GtEPTDNKzY5TFmlFmJk9FniqR09YpEHRFibDpxKOu3
7d+qiRb4Wk/eOVOr3z7ZM0WFCKoofb40IAXtF19KiqT8HtAIpLGkJOeGuDnu9md9U0SdqsrWg/US
Ie6C33PtfxDsjRG6Bro5qzdn5E4LCGVU8vOKKoXpfOmAAkBa1HDw7N3uD/8rLiN0OfB8A8L/Nim/
aqEH+wUVsTTfF+TB23I5/xyB+i3mZOetr74JNZf8vqo0fOK3sU3EnVNgcM/1wr9A20bf8ELparSZ
20TiW4CeA3aqzmaJ9MTdpS5SzQY4iB37DCNR6253fHki/bAPgSg498sgkeApGuXjblUR8aMmwAw2
0fa6GanuRCcYqjlEIhKYFCIj9rHqSXK5BmhXq3BSG5R3cILN1S22mP6kMITxrgNpKEzl9DRTaXdC
qU90VPddYNCPiT1bfNEqbIBxvo5lCKLkPtJv+Mkn1YGvAa3M6LU8GXaJ3Yuf3QOwHAnebsYJApIU
pNKjnBwHhxyOzudSTKaMu7V/nrQ54/I4GX2yaVwZmIyMWPyAaIBhQ5Z0Icq9ETT70bUX720ydiri
ASa7dfYatKwr/UjByIS1e9JJb8EFrnd5gm7qhpwvVb3GCyfTd4WKEuWMEHkQ26MzmdVaOmO1jfTY
V1BvmPWuTn6akd54XZadauTmo83EFcjsLFZKpeOh/cceEGs2/CUtFoSwfz2lRWx2N/g7PoSxAQ2U
6X3X2RRD3Kp8Tz1fbWLPSBLSbcd4oKFRfMSxKCf4gKNSnYbFsXV6EelyB/KaHgbBikQQRshixW+H
djgf1PMZIfM5kiGP2xYDmLgfdArC9u3IlF7xarEr9dQfeNMi8FNwqK/DnAetQA5X7yPO7ZbKzq5k
3rqxjd0KtEZmEZxp/XSU3uPGuBefKYyCArZfErwUcLyCc1ebHZVk3NMuxeQDlfgNT1IIjHq4Xrh7
nA9zkZ0cgTFDfq3L4YBLhSU5fBEoIyFgVOnIuc7RE8po7m6yjqb1Ih4jG/YgRhOPpqNlub4ECKBV
PcoNRFAGaXKM7vISSS4PSeQIVv7Kk3WSha3r7+9x9H949m3Ct0t2PFYBl2kXUWdU6V1biOLNZA2l
HS8e9pA+/g+c6JVXUaGmsKUa7Kt+GzOcPsluCn8/523viVmvPx6TCcmdiZOvkq0KJG0CykbuNVRu
5/xErPBC0oa8OfpgMfhdrUM34FsIsHnwDYU5EKosyNXgHHFs0E+kjXHwHwiAuloqW6hogcSrDZSc
J5zz+cqlVp8UmzpR9ZmQD7fK7euF2hS12SozLSD+QyJz7CdVWZ5MCBx6yq25qzDwk8dNzH+tsjdk
wd8ZeEjjhgJtddZUCoYd781HOTqgKNalhQxsjzZvF99RdoTHnEYl+1DM7DXKIspxGYDZQIT/5+cL
IL7wUd2YhuzZjGeRLuvkz3LhxJwSGYuzIB4kr+O/ZVlTHVp536oYI1NzMowUQirIdwUGUkmqOpIe
wkdb49GEcBmXeJoJAec3q82I/KEMgDUHSJK9SV63bumwfgP/KH/0Rh8yzmGh3CH1fDEGT+lX/yj5
Tw81szHVvCv8XBw6RnzbahNqvffY4+UinGrSvE4235K3Vdg1F17iyXHNEoJFivLqMeHXD2eyi90O
Xb4CZ6TnFh4lWjoEJmJmHtQyWQCafJnkRE/hiu3sLoBP9w+1fbY0rEkMQsisdmNO+R4EGu41gW5M
Adc+LucK0hqmfj+VdozWArQevuycv9Cg2i0jPusDzOb3xN10vD7qYCvfEKVQ39TTzgkEUfeNFqpW
3wanUGNEew0c1t7i4kLwTM1G1OzSoa9M/K/TZZ/duGOhpSYWrIsn9ysDYLq61EhsqXjF1UKzdvlm
MenpF1Y3RYivyLqlUbn+OhLgtJhm19xFpzA+WovpJmucTgMfh6bZudCG2iKAJLxPCF+3oUnerk6V
nI+J7Y8+luDiIPAWpE8tjfF01QQlyw+6WwSWJUIBpZ97/biOtJoigvztcUDMQ1u2AIRtMRQD+eX5
GYG1GxuhkKvk8bioGx5E1SMZOwMeZX1c6HDUzymaWi9sLtSJOx57CSJ74V82W3ykvvzx1JFmEFOB
xjs/OMXBFFCRxAZOkWJOhNzmXuXuqBmy0ooShhjXiNyYX63oL0lB3GnjrX6twLy03fbvd5InD9h0
ZmDc98gdDu3O6QqD5Xi5+JyLBJCjjZREO43/ZH6T9ONxc+RDSesvWzpEXECF+ko6PnqNK5Dq1xIy
BgqLBDPzj07jA0kfb6YB/Jk6CYMumuZLec8BQnrno9nM6TjlvPRDNmMAb1fKQGezDumh6Qn90FZb
Ta24/YWvd53WoJzJsapZwiKHGrpUZ+DiZo3S4J/ksmdRPKxtkYXIcUdokP2NzLLMBxa0RmNKx2or
ZeUE1194qItSIhngwf8faLgR86lsg9Yh5Yc+S35k3uOsknhmwV/SI/fN3EKoANSaAJhZ5bkAYGia
CQUv9xb1VcGueNtXu65WhEVo5IwHwlviZk+xt75svyloUr+4ULMJvqU05NJbxXDe58OCH2JJYVC2
vWrn+jOsP+gePb1ZiZ1LOYE7kBZskr+TemrF6y61dZHAK+WKg/k+V/MEYNzNzplvc9wJARBg+tgc
0n6rEcwgUCqfJiNv1LEf6Z0kge+XaWl1Nu3g+BU2ZA7dGXsDMk/rMd+LYdeZB4hxYjhQRKXFo3Ev
rLFWbvtsUufjE2CPE09V3ApWUzu2CKsshrLCnAmmX8JZZJ62J5sxlXMSSOvMPTPmIvZEnFa8Zpe2
vDEpj/OWgi2MYwzFfQMmc/vWC3EwpXtmqKpYo0n7zbOnRqdN3OSxB8mpCEpJuayDcvKTAxsMD+tn
I46+iBFmQeS+8h892UC7cv3StRFTctn+VjR1AetYQP57APbEBGB5d1FKLYt/FbUcwCTU/oJBmvRq
tXmHlsMRMeumCrsswkxLcbT5/Hr3+sSihPFFuJO5Ez8+BcqVq9CKTd4xjmtvMCdk759UkJZvMNOu
yNsIr0Iw+fAAW/AyF+LOersjfSRF0Q52VOb8Zvvk4TGBibiNAclI4ndhyVj9u/WgnIr1rk9/TLYz
/m9WfMwu3aK3P1ahmKsf6y4Oor+e7MsheqEIqIhicYjrq5Es5vkjS/lDaywL0T6zGB4fspbIIZrG
QP3XHokIcAQIvf8/gsi15CUcI7QbiONfn3aLVNXM/JrBhDBABHmk1NoaWIFFYjGfdNK0GByw0Opq
nNuu4R+BHvePWe5/YDY9LHHx0O8UE1ynyLeY1Yq0MPBMt4UAOM4DoI1ZZ90WFrCdCywaP8lb5lmo
BhoDu1mA4vxlOaAumXPPJKMShxIohTWQ1/Iwih1GTkxEl0Ij43IlAO4vKDItOvE5FE7HqAtY3wq+
rpvlyFN196EajloZ6fBktn5XN4E81+QRcBNQbYZoIJ1jISty7ZHDNOfUFovbRTWInNK3XtXvLXxz
nbMwjHSaDHXHnRTRc0mgceGyjfG408wC/u3YUrN6e+XxYeenRi3+i3VrkXTuRn+Ofv90W8qVGKHX
1wGFnk3Rqa0TM+zTpp8MOzsun1tTKbIoYYRGJ+X1hLa2rZqQD+KtZpXOz1iYHH3xsjFbTywuG2DP
tJFCDx8X1TO3suiYr6aS5m76x+xqqmwRBDgp0Lsb/R60oofazY06/hCGMuAw+d5hriNW5ur/8nb/
9aVcReTkjEsRI2kvbE4lXPP82OwGW0RdbFV4LEg/4iMBY8dRQ39IHn2gR92a7UJ1sStst8EamYDN
qeW1Yd6jcOaxco7VTdBZHQZzWPxhqUYtHXfh9c7bN+J4A2et0reIJHBaZEu/6137Mn40xxoN9jyY
eo/40wFxCzCsghkdGawWp120gzqBfI3IdGLS9jmuYV1Xeip0IoUuUSykJcnYow3C+lRfzpZM7g+U
y8Yc8MLhoB35XLNFAfnJ+mbEyRVWHleSISA4BOR54sUy0CEv/w+fEsk9KfJ/hEU4dNfGKAv7kKGX
82RZYW2DFsswyiSrkY0KleudYSpv97wHUipyCxPbdu76XNXksl6i9hcK8qjlAYgvcuADrsblHRpX
zRCC2DdCezHIeVGqjYt+HFFjqb4pA3yF4lb0AEnFUL2rAc5GCXy+yj0Xjiu0uJXW7NT/pVPlk9le
QeNE57JSTGkVFkVxl1a9g8g3tH5oETkGn0fI4BBk2I8c5KabQa1HqBQkbaF36k+fg4f88aDrLAI5
aCcFN4z4pzZtO06wcG3W3eY6Y80Iiiu4bltxxOQhgOh4j2ykqKUXiX4fc6JIfiV2x5CeZ9KRbefg
SAuDNdecJSCEt5iy8Xyhbigh3Ta+1Qa7B9wzVYsK58+8JelxYHmipHW9jWImjlRv8F6M6ZKKBnAZ
Po8br+urJSKTv8fObSGtaW2LIQao1QCXajW99ep+Tc6q1P6mUJw2GbQ+r2KemtbMz+NKzYfNmBBQ
zU906IXIEQRodRmJtZRoBnxLf4zS2IiHf28HAJDHp69gfQ3B2NZbmB+nC4LXsU9tNwcztTNp+ZhV
C/D3bPIzZtrapKK8ye2DoLu1PGXyx5kEKjfWOdZz/J7q2IwvC+eDnTvXcd4KwMe9kEYLpU3ADxLX
mWbx3hgY8yuE09ux4E6kSd5i3+avEJg9nCEDbYf2S37uWlGWcpSrwRKgBCt3pN6C0CddemzwldRm
YbbANKbYmHD9i0eh+GSyNQn8ldufPGfauY2ZIpOMQfWHiy728t0prRHpERO6jS2lPc0bc2uxJUvY
JMDQubddVGDDA7s6opAJ0TdmYV8ST231scp7/BZ4isUsDr86qb7CYsukofCPMO6bAu5XIzF4+K6u
1UGg1BWiAy5Km4vlaD6RPsRzlP8Pp0plsUasgwLXHCdRg9NiO0FCjW8jI+8Sv9/ebzwdmWpT3QGZ
PH6ukFBq4is/00rz3Fvn88XyhW/4wTJXbQ8u7XlR6L8J/Dd3LPTb0QYKzHVkCdEIe/9KAWTp6tJE
fhKl3m1CbcZeqstk+YVoqoxurDbYsPWPVSFsZ1br4/+unujaJiDEN4+0earLJUpiN/nM0GZefzEf
S4JFisuSXOzX4m7UuwBIVcsC320nvU/jCZmk5RJJegmMPtQYZ8QafBx6dStib8lgOmMfpfPdx9Ey
bo2bfmNJmAwZoXwUx4Uw2N89jKfHHpTi6VFkcFTcme8J81LI9Wn0TPNb4Ok/4kNQrCe7PVwNaru3
vm/EuZyjzI5YJekLsxlWTMUg04YeHTfd240R+tg0BHWK6Wa3e91dcuLfQnmIrKpu5nMUoDRBMYDr
BVghAN1YMalOqyoDXUC3gEiYgzH3qC7g0+iiUBFwc4RSLHeYZmq+/h49vSkFp2OojpufEINe9d+k
DaXilq4elb0KMI506uUBs/xsVXnvoNJSLCM8bHq7MmvGOm14Jm8OpwShPJ0rNcD9DrdJR/7XNC46
VME6bxjkgdx1mRQvM00c7y7F8cB06Pm3qpXdCGDCqXHctiX9L5JT5xezeZ+nhEKlSizyCmC5iDUf
AdUME65+q5X2vOmhi/FDhlHBIzEBmZ/57p3SHPcInTue+S2LZHKYfkYgK4DD9eatbGoLx2x1ow5i
985YUP3giPSf89+QpykymCpy9bERTysugAdFlaM22BWYlGM9fyZFmp6kiBZp/6wkfRTwbv5qaXIF
IBaWCD0Uyi3BvDCrB3pHsxkPW480aadAavmnxtlgY60njCkZ0YoWOsfP4rBeq/nxVhspVKtW5tDi
g8t9hC4Ma52POeUWhsrZGMazKu+WsSBdl8jomogYdO2g4EE0IrIRIbOkSb8flwQJFe7IZSmMiTEQ
staqZuq0mvWfDZbVs7eaps9J3nKdrWwqpZeLzQhlyAF2pdhARfey1VVay5F4/FawPtmNS1+Ep7uP
QCC5CHEL0jRJywsIgIGmCaqfjHUbJ4M/yojDkKcW7PHwzrK0eyRz5lZIWbQsA3Ystwjxta6m0zlm
xVjQRfXiXHv11/FbR9K0cYze0rzGuH/Egn7aHAWxRRJf9TO68jyks1M2GcBxcTQOkIftQ0NE5RHA
TbiMT/i0HmkirtHGalzEL2IwruZIN84P+3x8g6A8KjiE8V2bncZ0rWvtWvyzsLX0tD5KPSOaqSFx
50AT6z9A/V+YL62TmacrGJNfi7EiQtu6EmzQBgHUuMSiBLWgQ+NTIoacKex72lcvEl3wF958Gma4
a0cf8I9y311x8HxtuiXgJibx1parHmBRj834Kk2xkiEpbcS1oztR40ba6SqsZfIpC/GeXa93tw53
E/1MKegjl0FVw0fz6rmxGzo1X/XwPlkF80DSFRuXGgvbLxc6aIaF/SWegucv9zuqlvtm5WjkJTwy
m8Ayepacv94v9zovH3DyanpINEtEtn4hhfVexZmJV4AMdVyT+mwW0tHP2CrdYhFi5K4OBpCXOj2R
5oS/EnW7z7ssglu3S5JdpaIabUJSXBY5TOe4abVNavRZkDZpvovJkAQUF20MbnxaFgS2q4aPJyZ2
uljuDGcBOsY9oi3pRtdSuJL0SmhY4mY0LEEJevxKIRREIPfxyO//jbrwDtdZFxf/ng9nu9PvcvxZ
FB0yuIowLerip7F2Xvy0RWlq2Flqq3dNo4sCEg9z7lz4Rf7y0qFmA52hVqsPvnYf2rgRje+ntF9e
hHbL4zGmoWLzeQYZOY4F7fbG5LrJPI4ueHj74GvUPxbpu6haWbiLVHzby6HMLFHr94qoummBgbNT
7cITcqbF7/nyoIjFWPRU2t9bPSIfZ9kml0QlafoZhPhyv1lsdgtd8gkQQkMmt+9A+URXNqAzt8iW
Xo/DcR8cy5irolesnVwMlenKT3+SJdivKb29YJvJMmyL+fOjAA9bdVUcPkeSsHxotomFo2GHh/H6
jgJwnT5ueIUWPXC5GA4yyPS7eH6i46nfGtkScBWmI/pcFn58a+yYqw6NC7SMGhj23W8lYL7bEpV/
QM77KcU088iXL2DB5xNY3FAizhiAeHOctss23mudJGeldotAxPWqfeevGwgWpdHKXsuSW5GuZtqb
LUYM38X4Fg+wluOLbJRXzUtObKRH0HVTrKdJvPG3jm/6t0NM9pGGgTaGcgkrMTbTt3YyV6Col2o2
SB2OlhCUid08LKESV6ePF/RmNl7zCadI+pOV2VY9SoO4KQ+AdfnEtFCsnTxCGLTIctJn2P+RUrpL
MS9GPrDKEFLvXJClsbR1qL0EICVmqgWlwe4JweF9ErNtqgWDYm3HC/xD3Qrr49H5gqxkxIu9dmg6
33Rl9bRIcOSsCt1ro9o2IKA0/fXgSVwYuZwJ8AyFErn9/h3RCSBAMoBYAWSU1PmSuF3YgS9kj9t5
AFoQbWul/FAVxOUejYRwsI/rAaChQeLWzSrQmEsJYNsXOGBjSQPTXVeppMKHiwlYM8wo31kRR21J
1eOHivxo0GfKUJnv0l8q5+RKZho7A1SyUcorAYrxovrlqW1BLjV0csNZM8ewOoyezYOaPjeu4c1D
ypNRs/LNWSjnl6nQ39XPFT9WkH5QStn0V0nvnigl0Lb309sbPbub2QJc0uzAbutKZ0E7raxhv1H7
KZe54U8fhKwEopO0xSGo4VzU6TfRO8FXFhMwSsnV9zecLG0jlZ6cY03yX47AzdRXOi8SsgAiX/gN
RSAYeC2E9UMXkJOMMXChIzvVbDJPm/sw0b6QTxv6sY5sZjfNt3jrAmARULs4tyCJ1h8DocmvVMTM
IR25QsD5SvPiCz6QG9U9Ks8MFRbdSrWVsslxUgD9LjNRWloDsVIXI8S/IkHZPA8MOuf4PlFK7qiS
fWLgPRcd1AUjVEF9/bFOG5OLzSwlQrIUnIaufzj/d7EvvIUXetbfnl+7/87OmSjrwiy4wtEuHsey
aC5Po7NaL60TTA51NIcOxpMi9g7fDAlp8OJdOm2HMVJWYiGGtx51z7e2HHSqqyoXd2WXfp0hXeiU
MamkaPSpK6Z3Nbuk+nloOfVhnnPbK6XoELPMhHQPcDANyz/ObYmkNb9hJgILQK3pJmSbDdENpKlv
AzRcAnxGyHlg6372Ax2wZ3mjucApEZStFi7Vb9na937Bt83/j4/sdvh4HPhsy4VEHX1ZDmUO7jLI
NtjRynnGVWUjoVd8BRxkmpjBtikkk54r5yB1FAfRcyQTCsHSZHHZQjqaLU8FvJHWiU7aufFhqdyE
a3KNhzVC/KIeLk/cuI3mwPkrv/CuH3vnzwPqrv4C7XsEK3Bu+MoCjVO+b3hd7P7PE6CovH/ecYNq
vLw+05uuuUZslUdpaSmPpzqSUb9ZbW06hLYvIuPz1evH6oDw+acb5VTAgKbBh1ZRjHuo463/Sv5A
WnIy+8cH3/hZyEBT5h6RXPxtmrHtvELuy3seWG9O2Vwi3rEJTa/x+FEJfvJ7RsiEnlESmXucTpYZ
GssGezNz8lf6uC6KnbgyjZo09ToaOM4vnZbgLdjvV8ur3XonGOuHNDo06TjDWQgAfVmAp8G0tPv5
fPraBWu7599uh+QG4+2qYQcplz/L1mYId/cGFDjFiCLGG+4mAHP+81LRn183G6S36wzM3PUYussu
l8bhKkBp0MkZzhpnLCClzYLZ0J6koWJpJUB8aBh8IIC+9vEVzi/NIaWUdZl4h0jXPP1yYz0kdWAm
jaCfPp9ee9JX7du7/NHSUkdIKGNqeWQ5Ft69cz/5JxOt8a5us0xanRef1rXxmgJuEqsTh/SsEsaD
XIW1y7caBWIiE7ZFX4WHrf34TRoXbTS25Ft/1WkIucZ+BvZ4EWq8ZzLOYwWlfs78cjYyNLVClZBp
uiDYtfboYFib8P86gSCjOoUP9KcroF8byVFRW3e4NkkXKwTgVFOwN7ettTTHPBRWO4sUZ0e/8h05
dcPONnoKMwhozytXnxi5hWEETFMDVuA7aJ68zoSWgLYimrY/A+FlcGxSVDXWb4vWYrQO9ACYRvtj
HQnRzkea/KdKsa30b7v1w/9LHKlmaxTcVir+a/nguLWQMkYQ6VXtUvVFRRcOZnbPATwZWPRm3nHb
iShW7oCjMe2t+z9XCOgTFreDij3v8rFsvipYT4V7njky5Fe2u6ean1RFMes4VrlOHwXc69sri0UT
Z+ZFtrUoJJP3xkmR5Cr22//VXZaIsJr0SA5Cs+d93PR+YrC5jUFQ5WP+q6kSVctxZvRRJgkKZLRs
Ix5Kwi95WXAmXPnj9gkWDhEDJcAsyxyyzZw5L5S3losMoqMFz3vWfeUHskUY4xh2xz2hkDa+6Nb3
tLKhIxPQIdK+CwitTSd+KOZggqArPiBsyZibuA5/RvjUvIwng5X0kVnHNhhRKRhZirfrC0L2INg1
PzA4yihmTwZlb/1WItTW6ipVWDTRsfeWuPnCym5cQbOQ3ue5GWovKWxHfdJ8qvYJs71dR2fb85aN
k/awmSN0nBqnQ9AiNjhx1umnCKSD0t0sCuynH1tKUMeBmChnveOwNZkT3R7WN3KaXGNcwczftqJF
6J34F37+beJxp/ZtgMp8mAzXp7r69u9BABmhRlxHjssQMj/MCLbffI3p4wnKk05hxAM5JWHepuUM
D3KcIJV4z89CEEJ5YbNH6oanYZ9ZBectEWk6fWIE6EpDEDETagBL35/sfLS/MhbaKaKpLt59Sc82
F6C4M+FCy0LQV1U68MGiO+PScPfryR1a3sratIEolekAmTRVobEddvNixlVNXsHqAc73lsIELoqf
CTPXKrVhTMrFKqlytlxG6awLUZu1RF+tRIleWo2Ub/d8wQ9gfUi53FLmeYCFgGEXDWwtdnDisdmr
lK7vMNhhy4T1lGeS1Ss//eRdYCMZIEmj9U+ndkPJKRCzGDk4XBYL7aRTQr0TedmaAUz2dz/ONSHy
K3HPJHAvhpOaSJjqHR1pO+CEzbbXY6e/y8FrcsYYq6OE4XBSukfrOSgVgOx57nds8kSjiH0YfNgv
IRP3F15BLCq6G9Ytz9AUvcd02qfHi9lr6i7gIBS8Ml5wthLXGddU3CqV/aPF1Kew8FnqLSWiA9Ju
N5zUz/nO9SFNa/cqeTFGs5JE2kByszp+V25Gan/4fFBCq2cbFozhWI9wXt/Q02kmorYg+WlUCNZK
5m2k245pEKJ8dWquRBdgM4Nd2q6gPGyxOJ10rBEFV75Zdkf9MZZJHFFRgfvfc2KCLuIbaPWtcXy/
zQsbuN9wznTgghRUEYUJckewFkF7G9aOmI5Vc4kaSjvSI8s5XQA452LSbJpBXfzszv9GKlpoqRZ4
kGjuvCidXjwJ5OwfdA0aAz7dCei9DqpQVj2jLBXBr4C4gb6lXOD0EJSBM82dfDhXJNTUhH1YibEd
Vtylfe8WyH36BNVrL9tyoJlSrh+6VcyeBJaTUtboOzO7ExCaXcSJXiwBem9RhHuwwhHFFvU/KQlb
qs2Q+VtOkNo3vbtxxF4izK8H+P8+uaINYOsqXHf3BDFaSH+V+67v0+oQuV7FXtoD7V7QpX5nJzwU
LFUIA2MZKOf0xsi9UHPiQDgoNlG1wHFiIysqz8oJrL5NUomHE683HwsDHuJ+kvbiMfiaV+i9cgI1
0i5A83nTRVLCUiL4uVONASS3+zMKusbjixWMCUcNzfuQ8VeOVHX3lbThGZTyuTIhgWxCfa0FT6aj
Zqs2GeZej2XAh38RhOL+h8VBixZkAwh3iHvddJjGf3P4lDGTj5l31CQSYsumRXx0LyMfeAlBOCxF
OoeVSG7TaMsfKPz3DRqA92NszH3nEpnPXvsE5yuM8fWf98FLgNLaBJhP3VzM11uC2nkiB7x5QQeg
l7VESi5AgWnbytNpyBn1mgdNH/z/JVZWLZlNyAFUjC5a4E4i9Txw/qa+rDwcxH1VSmrGDF3HTxhD
VkK6rF4GKR9XetC4KZVr1fStEVAuO+E0vz8+8N0g3gqwojRz3gbEQ8MUhQxKQR+MRpvpc/aK5Rd7
GPTezh9nZKaLGimns4f5cKlHEcJDHVWE+8Ll0VqSo73IzR9ddoukXDDOhB8wLa2GWeuI+EeKaQXq
pw1xkPfZmbXh8hP8RZ0TypTxL4xrcZC5PRcl/Gz6Tw0U+86zfXCFRK4LLNoTJz2cSdbObkk1XTku
rRIOW2Z0AH8USc/2Vx2/A+zsj6V/l57q4Sjwsmqz3zjIvLB7kUMMp1Zth5ZUo88a7JeIrg6Jjie9
Ew5zR41e8ltKjGw6f2pLu810qjEscSkIz6yWFHc6I40aoMjQn+VuFw2SdCuw3rgA94Zb66PXzbgh
tMNxtZKI/ljFMQdxlSJ1Ua4omh2SSqq2d/s4inEup1RJu/NCnmo8AgUBJPg0x04uEWbSx+tp/a2u
AEhf3Xzf3iIp9XG4ftLQWl1cT/ZpG9bDczcZuyhHHVBOw5y42s6oa7tdzlRRGuT58s+975cTj/JR
wUIK1ti6zP2gc8i0BbO5cG/iDV4+WISHC139Sg8v1JSPmeVGp0777HWQVbrJVDoKhBnHYGhapyg2
c+4rOW9CrAI9bhUJKIYOQk5/sq2fljJScbROu+KahClsd/SzmCaH6Kx0VJSJPwxaK+yv5hDtSIZ0
Saq4PU2OSdl8F35c1iAAeYg6GNW7FMArEq9DtQvJVNFwFTYqC6Na4rj7ZIHrRmA+1RrFWcavLMlX
0KyXEleAoGZE+X0uHp56xiGGh6PNLnDJiKvZtd4fW2OCKjZmPgISxcsLmgIINrPdcxidrjZRgN6E
dDQe/vyG9J3D1P+nehRgvAp1nGZl/LL1rBMjuXf5E5soHflzhan5WacGCuTXmBpZ+S6SH38pbi0a
xlI1h1NvkbhOuLbBgGfzMNeZgqtlGAmZE/TIRbAHYWXWGovU4UwKLANYc5vhK/eeMFoHO0LtjkJG
jHAJ7B9v6hxLFl1Pa9cIm4rfX5iM4N4CpVSo6YctiS1LsprucKb6EkeBmbPPyV9X9GGRwjvi5Iad
0O1+WLWsc0QhkUSpqVtA123G9MMUz/GyoZo8bmyG77YMKlKZYuNpgq6W/Kvszw5osDj2jASDmrxJ
j0I6pkW4lvVT9wo5Bo2WM7/EvPXCaHh/mVRrI/bpTaXm2s2KGHaXZq8YWWqfuyLcG0tmD7o16ThN
/2ocJebuSC27OQV8e2g7tRihzWZ3g5TXO4jzCTXBYneEl9JsWeeWXYAOWQ2o+LV4DUt2gvqRcXg3
as175hjpnRao/R4j6C6JlJMMyCflgRErxAQyydSXYlkOXf53GZ/DLepx9NIJjQBLbyKWQtzc5aXG
wNpYb1d61mZO79JpTt3dtUAF3O59ZIW8fTZ3Le4wb9Skepx9/LpWbQsM2LEwhGOnUYwBIYA+aFHJ
TZGpFUKHsNizz8gkygc/YgW3iiyVH1vsFW+NXmbP9rjCMAqQasMO/rIJzG8w8hDdoF0eS6AYZbwb
pEyNSvXwSj+U7GJyRxAUcnf5g8r0gusBcdYmKUv5sk29qpB/4Q9/mbrCKwjojy52xoKeUmNYNh8j
Bq3CGgpzuaA2NtOSlsgjrzRofcQLR33ZDRKqnGIunL/zFYtZviCV4m0VV2SORUUJaXK3HzSVqE/j
06HwczHfORb9UzfqOirjOeg6RcfdsntmRPNjT+cDNBRXSpYr5wcPsSrp2H4AcgLQL8QvXA/2SIzL
li7lnKfa9O1AFrdPG15ZchUU5UfgQ6E1vdIY94/1YpXSKeIOwxEhIgCpTb3qukR6TjFLjaJN9J4Z
KhzcjWI51yWjHTe9j8ERhZGq8I+XxJI9zmdllEhu98qEMg9MA7/e1PrVyq05G9hnMRteDFR1cRQJ
xFbbblPOfbpewfdH+7BRO3UQhdS+hdZQFEzk1Txpp3Bmc3LoW7bj/QtVW3N5K4573sl0zHWz125P
VRXxwgP6L/LoNuP7v8bwd/rDruytBSpVoTtjhpiuQMQryk/BC0UFuS6UMqFVC/tmA/M2eAgkRHES
fTou7zGi/7HtRWb4wYW4GA7MpcWPtN9ZTxu3w8LMPO4dBSlmoRd5xYEn1D7cJ3MYHaXWrDX0TtUg
dQpj9mC/d1dLoNOqLz8fa0Q6wcxITJX380buLegkpgT+E4K+ZuiDZyMQL/NLLEBNRPlw3sLHF+Aq
DGYiPSFg+8Cy9CkZKBXtB+abkP3Wab3O9rD6am8XqZZ3Aw51OgZeglKYtJtvZiD6nDPM5iHKs0Iw
3a7XMlTlo1Ki1/tuZgYHqCYwdbKtrVQy67hvydEeE8FKjARRa2HQcXV0vJDlIdPNoHnWaActgiHD
+QUNcaMl6v8Z9Aouqms2mpFfJ9CWr2hc6PSq3RrkutJqfaL/qG7CQMc5Pev52CYSP/4CrN34RKoI
PJKa+6zpyzvGsBeVk4VI7HKPyEEeUllznIY3WImmuzIlrfuizLdghsx+zEZYaofIYrDeVHJLamzb
dmUCcn0nKeNMqr7ZLNxVTPFeB6kKbSSVAsaKB75vhb4iYlN0sMoCF/OSwV56evsWXFcATv6sEBUI
hreKr5ZDmrN5TLyi8g2CwgB15C5TLsecA10foV4eQnhGoxUvZHehHuEGdY3rAaMensR7fCL6ndXX
QznwyRksFR7GyhUYlMFX5zNuEjBYAmlBcDt6tlOHBCfg9Ur1gKTljkjTbEO/xErRvcCZk24CAEOn
xP9pSAIdA4ocXYLQhBRwoH/0dgwUAWfTm7B8lwmJ8mEOGQJ+AmMWufstP5PWF8s9E7OqKgCVoHUY
fGIf1fNaZR569hJoDY/mXMQ2jVawJ762FtIPfCjmWdygBf/EhcUkaMCvzbfRkRqkCRzaklnvWpba
9oG9ZPnqMrB7RXaI+gVmdcEjanwrAwZ7Qjsh4CRwCquamKXZjhYR0N2BM2hSHYiHdM2KJsTQE9Lh
OxfcZRGoZEz17xo+3xyj0DqlW+RYfYMQdPR2ickhcc4xdhk45z6nvndX9g02nWsCg+YXpMSYAl8a
ckuEbkTpBcMuhlcqe+cNQkF6RoGeEsyHKaPrBnHQj3hjelN83BQVEz5OPBQMPp3m4iU1cOU4Rjc6
SSa2cuKipU0dT9CYWiKhT1drblywsThlpCK70xBtD3BA8EbGGW1uKkBNI/n4IhH21tBKiiVQOqjN
lP2Uq/Z5HcWa7W++w+Mxs1i2o+nGc9ycpjmRaFjbQ58QTThMfNl1pt+QQ+hIl3vdZRQ8W/37M22V
bopOGa2e5wkbNavzlA1SXMsmDXKmeYpa+pG5Pk8HgPLgsUXcGox4RkoZa7uVlBb0PNzTFvjRsVjt
fUnrp/+d6MYYIOuZfrur0VnA+BTntRNZPPD9tb1hZJXP4Dpo8zyGmBL5zo+pnxHqkwDwflHs8qZB
zt36ppHDqodyLDgcDVzezyLSDNRHyhI6Use6dQYCNoR5xJrJCqVmApugLlosn5Prs5xdPI6VZuIz
NyGCn6DVpd3Ws1p1VxNJCW3a2+euABM0LfWWZrllLl5QVHLY7UetU2Nkhasp/dQWqM3g70bVTMnA
lUKkx5LGPtyKVFvbGYIwChbwW2Oy8Zdt+AqY++OF3iIR2hG20Vq4LzxtJn9lXM0iG13XpIUgN2ZC
pU244n1T3JxwP9T2EFDID++eeVFmLIBK0NpDI+m8fC+8T9WEArMxn5FKW2s2Rg3BE8irqN5Xrb3Z
w7LKbw8jABK5c6mWPYLV8R5abIIFwPmPWyRU0siFzcMvu2IrjQ9ZCpXgSoeXduQCLpQKzfpPUL8h
GoxPxn6WFT/8NKLTX+ECEXFIDGlxkRRwTwGjAGy42BCLokw8KW1xGX2LQBEweTp7I3N8VRv3T9E1
a86EWcj+CRIEgxhhcT46io0LmaHLd8U1jkyi2650uLE/uqwBMNSmtcmFEC/RZ4RijCKSGtDbvbHu
mro5lg9YTNtCyeZ0sGGHRy5aR0tNV0Ag7zAvlJG6cSkrNrJvDPeoLKNabpq0/Ovltsdi9rtKtKf4
l/ocU7T8xpMv+rGwKcqP2glF46+39lTNeKnrrCOLnyBmBc58Gpq8OihCGfszKIdENGCdMATY5Ucv
27x9DU+sE6Npv6ZglITvy9Y5PQGO8I+hua2a02ElVVuRl/CDMs1SdQvNdb7W+jMW+s2AAKZweu20
0WNe6qyxJ/ZZhdlKgPnN/tHYvBw1EWBvfU9S7vTUgK/TY0Sg70kLP7dS1EVEbHYYR3kCbXz+piFN
CiySPfSpVsTl3nPoINpv0vc8DfPnAC3Tn8rNUHw5ynlrYu5IGWKxhtP410EaBcLZD8W6l0graEQD
Z0c0VHYC3D+H7IzB8Pvsw8BT+TinrfXXwAxxVoRZP4fEcLNjfQbNr7aGqc0eo18oi7XLOcIVn1pU
fry6dW7V6ecKCBYrbyB0Hwn7fNzOJwhWJmUMhhNRbY9VvuLaLIgCxignwMOdu2s1BDjCzBknVXce
1i2fFKhN5DldO2b1UcOSlSD58OCHDqXvt7bKq4thGAkBZa9ECi8JxYkFcVSckdmSBgpaeryf0c6l
Cz4iZ9J0lJD8D67M9T+h6nwqu+0Fz5DFzS1pzwtS/1w531a36rc7VME8u/q1ohnUmmM8Hz+z0twu
ml92YbybBnsFw1SHF+S7j7dc4Jz/0G492qZ3lUkSd5GbVGTJAfvyXYcFjCVflTclWI3ZzK81YWKX
Jh1ZUVdR9LDp1PXT9AVEyOVYHn0YDdadiTjz7rlTH+cYeYS8iqKKisMGIGuyaSpk94/Euy491wu7
0GsXnGArska76y8JG1bsfaoZ8MebhGTwgmYUWblriSTOtqhmAM5DSygL0V5GkuoC7+PYlwCNt755
Za1Q+fFNqFkz92BkCSlnjuon5B00syx9tozMTfglZ3CaMhDOQz5UfUNDqbdTzbLy8QPcxyfFzVh8
EhlNftYYW1/IjEbr/olcOHuTMaQ3JJIYPJzeS7cWDQvUnmwrKTL9lKedGm147AZwWJpy7X8hbb7C
7VPavwPF7W/4dcPXVsHTGd1vqg16S0CCA2j3csgwewA5aF6uTeW6DkjSWzaMglxVAtKZuxQuwFzA
y0p2E7MXBrctB0oVmVkLCku3ko33F8Kp0UcUt+loYZfTjvFP5hvz2KvE/BO3Zc5HutNptcBkhWBT
wSAu/XE+PW0j7uqZeShVdDD1unir58BtKKj4paiEyZnKoDxiiGqB8srP/iNTrJ/imP4cZjRRGcpP
SSORJaukYkfBXC3kYdZA925rQTyn9jPeTi6zvEStHEb+kW40XdobAhCe7WJ74Sl8u5RrhKPZyzkS
1rNW4f6O3FhvVLwyT5N/ADVXAoGsN4ceHwtxixErmzuG0g+5c9pTCi562f5COv9Dah0YP+86BgZy
fMpq4R37bSVMJvHCs57lAnHIokTzdxcQMSwvudkXda6+cq4G+EmcHMXTlgO3PFMtSFZg1LvYQzoo
s0bnj0lQp7/yeToBj3EHXKbLEt60KsS5uI1/rn3dc3diwJVvpQZRzaU5I0Cu9nSk6tTEqmAso9Z5
PsYLGBdHg1CP0bMXbwhEWjf36gHCe0/BHuNkUeOHDwDUQ2DS1+SHn7WsVcCt2dLy8mvPBJgwzBPz
s7TRleZCONA2pbX8gV+bxhZFLwO+vA77fA87O5mi0BFvTP3gJ7LIlAPntZ9jd8NOMJaJclj2voon
qx7Bpsh7d/TV12W/qZe8rJZy1ZW5tu2gvzZDjQ9vcWgm93v2liHwFCcMm4VN8uyCOmM3SBjC/VXK
igPdsGtWUje3r1spLde3Z2grhaQVZ4J/xCPZX8q2XMkACs5geaoxAT2qq2yI1VWUGR69vHOIuKmW
8JZCtJeU213bPiDk+CyREpY9xLFvVOYViZhdFQPbJOPAxv82gImuElmEosgyK+KbpVrXgDvkT6tw
3oGxeX29ZzX+Dg9fJHZyRHTn39EjbSsA3XSAOscEFJXS3S03T6qJZ4jelrQ6NAg7sKJoKE0XhenW
rxSQGqW8Nm8kzR0lRMIib+VBQse4RLAXQXCQKeC8GD9Na4boqYWtV3zXyp1IpVUkROj03JyY9552
HoSkZfxQhv9sXU8QCghjcOzxMdcFJ2AIL1f+uMilE1D+bCPV0JISxmp+VuX5mrR1LwVDdOcaP8BW
ewFoNunCh6z43L+FhjD9vMVlLKvFvL9SFj2MMEErb/gIJUzALvXM6bYW4qmBMQN9kJUwf0MpcbIl
wGovZxHfkq+cjtGoZvBsvSnOS1ep6y6/hCs8LGgfP7kgbEJKFrjMKMyggniJ+v1NkIArK2IhL/Wm
Rc4hZX7cJx7ySLml4Vj0HprLcJZJHnzL8FUELJXIl6AmVMq0t2v9w77XEYcpqvnPZ2+DICtuPJsP
YX+NBAQIoRTgqho/KJDbjPHX5JGSzagnvCVgHoyEfsyrCYG2qDJlAJh+GVqdBztJLcnrQMWEpBPk
3icKJyVrGowRt7EQlxALCr5Ze/+wIYOyOaYBVQKyyiIIf1fLEX8woECBVEv+RhTPw7gV/LQgjTj4
3C0VgIBpt4JOboJXEp8wAYwRz4bKJuD2JLUdVITqlHspp6QS1/Xsawl0CKX02hiMrq+sNeRXyoxo
7C6MNCaMFJ8GyADojhU5B+nuYmldeb1dDv/D0Dij2vqPHMRI5maKH1nZ0QxGZCyhMnykvIaV05Ry
tZM0gSTBSmhG1cLokE6aQn5/a5P0i0i2GyMwulJEG08vl4qBAX7r7/KSxa4OJAOd1GzYWOnt2Q8P
IMcpGAAsK1uOkxiw/ahIElAMgn9ZPwvzGFykECctdwUyigFW8Zna1hHjh1XQEg7JjfizIMzt7JcB
vT9CwOVREUeHHi7mMqtrKglolkpFDk1hQO0PTrzJbfGj0q5Eq4sP66ZnRH1g5mVGR3onYcWejG3q
41yyIO+YRrB0gusqRXPxvEhg82AXesFj/Hrl1sm6EXCUnQIelyi9uahHKqUwbyTtA9+v+VpfRc3f
wVuCstEqDdrSqT24fmby/Ys+XNvmcjU1mQu6/4BIUbBi/0qcAaZTVtXkIHs6EqMg8ij+9H14ZHVn
jz/e9ktc+GZwW58ZWfIW5cvtDarKP+Lw5hIBfNb5Sn6HurXHSQK32EXMW3BEbBMTBdUXsI5yOW2z
CJgqZ91ou0MQOK5iZ0UO4FFUPejqQFe7o7sSIzdoV+OS99Y1nDI6bg5sUeRm4BiIje8O0E0mx0Ru
8yjbrNDAreyY3qFEvGWlnH+CD0YkBpnW21ovUU576QDUw6+WYp2bAUKNP9CGS6aAILAcL7H9fHi2
UaWcquaafEtmd+8Xi23OFZleoNvjL+QAxFMldy8bU38mhFiPolO85/3V6dqDKit/nIEI76xFhDHd
FskCFFnZIsizkwd1+jOHjKbuIxyT1JGq/fkPH8f3kC2feiguz01fLHWDtB2mo/2fSwap5UPSZ53E
u5Pcthp/2K+JBz10x2pJxUVdiYvzgXVxHJF5PyLoOA8CItZ4Zrb2evXyrZMy0HvZJLYyVKKkcjPU
gHsIOE49zjyLiIejvVdT3LDnxW9FhmvWlECtzwEku/6k6UPIO90UTtZn/ACdIkP/WAhhTrA3NlG+
9OYP+f+9e8G2CUDkiHSsrxXsowOmEAYxEKXcEJA4Ch2N1yxnJEmVxLVCNyXw6Mh2T9sC6AACkE50
20lVPwfl3AzxhIf9HBKC2PoJSt0Lqpix176AkWYsXo2PVqplEaK0gdVPx3SwnSvoA+0CgLuEhxKh
VLnHNlaaFd9zohFizONcjfXvTyvBMl25D12XSZxYuR9ovPJZ0V1kurPH8crsOCn2cHtMaNsfllSH
rU2dJoadyocqT39h/VrOwoPuyK5lzwAoQGTj3+l7gnrCyLQ/0ys37VMVRv1/ThkOc0ZETM4tdSkg
RhZ6fuIUO7BTymdlv5x4Jn7Xbq6SXrAe9Gut+u6/0dayXF0trBBHSFXOkvHFK7E6p2gcJsaKGRd8
K6xEv+KJYRiahz0ZsKMtxeN+PIdDxsqy1NZ1oAtRGuQeih1zXSUDGInHY9KissPZoKct2WuN+PHo
XZNSQvnri6S+mfcXzeREw0fw9YFKNMsNWsUu6Tkm+N1kOz8Oywe+VORQqsfEdrI+sY4Y/nRMql30
eMc+4yP2sV1x01GCSabrisUlA4LmoCICweZXlEjSDXktjg1v9Hv68of5V+Z4WUrYS6qDnxihAeNn
d0C98aNaElUfs5cAMq1M0xDOlvc3EgUSYSAKYaHBzqHOAzlFgaN/ZCHPK73Y0ebDMcnHoAtr2MRj
5Rim3ztBFlWgM+WAJddAPN/rw868AL6sJX3Or8mjJ4M1fKkWPywjrEVNosIhUNls8F2k28+MLsBy
Jw2umSggfkdYwpyrZIhgEPxQWZYHHl+9Jgh+zb4FfIAwtIiiTU+7bMNmCUh8gX7hG019m8XLXaSN
GbPz0AburAo5wI7agraH2D4Cu8fOIkaAvKdgTRq365cNVTouMDiIpujklmkVRH6YPT5hUcCecDqZ
Ltg2ZldRb8v9qlmYlfxGaIaMRQrCHQIyRj0iCl3KEnr+Z3XXzzCqRKjqFmew2juMY6rgPx+KHlz7
oKDNQzpn0UDZOpu1uavErvoIjZe6dZ2xErtXUHxTf+d1F0bf39SykgPszV+w98XtuRCdyOprB6OA
ExTo93MfLgNvpZmTXpGy4xFPBkIgmYj5mnm21nDRZwQvsty7VXEmhwTCx4ID7T7WMr68UgfBKVuG
wugn4nrFWOuGlXlmstCsmmjf+0RjG7fpvOvZ4vlNQntbwaC2xhWuznwkYMM/l/+imDl4fUPnqs4S
Onrfxm0kg06pgkeIACQjCPdwt5NJI118ytPbpDGfHbjt+A2RWKe+8XjlvLJTePhV0xI9qwZCM32k
tUz0N5oWShq0s/t/kziVuX9zfZwO9tRuqhR339SR6TRnHDUTx2cNDQbStAkO+w2tMy+1PXKoj3py
77RegO0YZmmNrHFN7tBiLY/Uq5x2RMda9wspoOwI83S9eQfZNloM2XiB2MH0uXtSJrqixe5c0NZb
SDIHh/IRTuoM8d9z6mI9ZzZoITlhraA+47qkAJunl+S+K9CEmyHpwWr/jlX8r+JNEVZVP6GHX/Yu
t/l5ysc1EX85Q/40bl9WSQQOmcBytr9g9os/nmflYgKLd9614BF4PNE17SKgV5+f8xNjEL2z1MPX
ifT8QqtOe8n79yVYvwE0AV/LL7Fztpjae53WaL6culL0rWeO7Yty0y7jSa/X7JbpKVNgqweDlWNf
QmbcqGhj4fE7opIO2rDER5VzbmWynXGAn6qVhTEbOWw7+H7rCsjiAaV5GagiWqyXxIJaXq0INTLM
fHlLZZzDtkDdQOch9cYkwhKDH9MWksJIxCTWoSlag86IunvGRCzd1DmHcDw/RaNzSPIaxYkPi6FF
cGf8DtzpwnHGp0Lw4KSCEQ9c7hsw5LzHx5dlEXlKffmmwImMvHF3+0k0biAqwCqkJiNvNKy+fg3o
li5zMExCLElM79nN68wt2ux8vOdqxJMBjvDgPeqM/bYy8mOGb7cDUMbNAl7gWvawkH03E4l0mKxE
nSugKC0HLn38v7vbDYhbkexfhOnsT+awzmJ6NvPUWEOR/0sWcNGSIm4SAMWPJEKijET0Mi+6RWLP
7X55SfaCKSEfaYHLKsdTzfpy1rQq9z5MLWI5vYIcNsl2TGq+truOByvZAPSt7NNdLogYmemnvDgS
Pahr8H7km1sGfDeppHGf+uQLG0Yynzhx1oKUdbTpkiYIWksH1y4pExLeE5UhRBhNLo5tJt7LL2rP
G+NKD8LwYvXWLwtnxjBtuf580EqjJ2blSNIFGte6KI1Q44sOLy2vZ7bLqQ/w/LLtuM+CpjGc84q6
su1dKEO5UbeVU8BvpLAZ5qLqCDA8gW+GpfQP8Cj4Udt79osoe6lj2STr8IG+4lQAvAcAkhD9M5KW
/uc94LPjUP8HGfmuD8L2v1sZ/ziRl917lBpaTU+awiHP3vxslr61XBRYpmMwWHQTy1YvnKqB79s4
tUeRqGikf7vmjzxgRXE0l57Hxqi7GrKmHjs6iAEkCVshi/MKKQpdzJ11Du8iRDfEZKnTVHYY38QC
od8JF8v6C/ryY64VhggmhnPKKeD3YIXY1j6LCjOXcUbwqiItkpHwT/E8O/L340IX0LISeSqXNv1q
i/wvJMm1JOxxuJZ5aLnBHzP0zpCC4o3b1BOl0YhWJMA9V4wi99g6c0jySchgIaHXn6tV/Vuw6lYH
N/RL/VVMYaOfO04BmVNNFLJI04N2S7JceR62JoE+lvkUPZz7XJnA0gycttR3IQh4YYFUctoiGCsO
llGM9Bo9cZpeT5r9NP/PKsGApQC+Jk9IDKuDwnu628GANvDN5BSok+pcF7TNx4j1Ksv/tWfB0Pla
C/wg0bDhAFOJyE1Rwd4Bc7w08AQOY2dV0dj3nDKTj4BRSeonFBLvTzE5koSvbRsK1DV1iiiLOztU
GRysZ4xCILiXLCpRsw3mIgqZlQU2v710BZ+US1+7e9UMkzRo5fqiZrt2qZgwmuzVv/fHN6iJkMT8
5x+ceAuxOdkQk6GVR2GAVRxVue7hj6jwMO6JXhGN17PI2FTI2/nDLsHefLsb0cF6qgLNIF10rxbg
vs9yWRXLYGEYqj2t9x2GaD6yZAxGJJTj5RRRYbBrVUAFT/qNtI74O946GVHV9SFuAEQzn9+LxUOc
+KDG5Gqc7AitNdv1EOARkqrlc/AwMsOLkpG+3YBSJEiaOutMUCDhqztCrz4pFTp78ZLIudvyHxGs
vT0IyvJi/psNs17fvn6PIHvBYFm5vA5NiCrbi8J7xgcNMNDx2YSmXHVan/BH9AozJoICpk5McDXs
BGIfnE0XNJnygV0vdbycrfTpmdVJQA3F5OyXN3Up+YyypzFvKcpNVkyaK+I8Pff8uNV1I45dY0ZW
bnqsJj1pc2JN/Mds9MLYzMyh48eVcLqz4s69cPYTgZA90VIiHATQ8SAFRIvWj3vGJPg6xuuY2gVT
7Bv7JM5mn0quF36CJiaa0qMrtvnbEHYfMJQhK0o3TScpjSBcRHU80jbKpYwSXPOZ/dSdq3tk3fEI
twUimDcSDEsC4wkkCuxBRcudfBV1+ahzcyq0Oh6eyw2jOXIK0Ea/+/dhYPASbG3LpsUTFjnDWHPk
POAmundowC6lneQAiz9sK/kEvy7mvSCWiqWpWLP7GITTYawGgglNfw6h2d66tV+ajLteCUitXBUS
MTVQc4x4pvMgsl48Akc+Xqbn+SSbuZnUoNs20uGC4mDIzPds9mGENWboaTimAxiy5B/g7Faqq7vb
tS8CkhPSClmHVk53gpjQ9hSuyi+ug0a6YKyO25razMsBadimE/TBy/bI5JA/SrLF/Ff4UA2qicnL
LNtFnjktA7kgJsayUjaiIATBGwO8LJbvFS4vkWqg4xmEGCm/HxDFYk9/oWwO/A/GHywojD0Na80Y
/8RWppCgp91yNyqHxfCup06VM3Z8syoD4LE0GkpaiQOF/NJZddCGApmoOXh9f5HN3oIk4m0JDFio
hHiA0DYhxhuh4eMiuCoFVdS5H/Cq45L9km2p6zlrzbZD6wOWP47YFCwwDXZq8lu+Rh5O4EA24not
r6SNIZrU2gBajly5xHro+9VGrI2FN/rFxn61Hi+9fvdJP6F9iAh/uJPf1kY4nqNiQnP+9eI7ltc0
c6Twi6xnzbC49Pppp2yUbXt9sLyfQ1WLtsUJpXvtVufBLjsQn39Glx1TuCdx/sHuA4zYc+assl4p
G5ylc7mMUwiceCNbLzg+ZSxM3NIu9nvUPd5q7tNMl9FZrKgBHyV1GBBVphv9KDX0FvVTpLEPyrmB
d+Gt++bRj3bEgCwSnOGZjFW0QWTLmd9eBTcIg3MBEpQXqtwnRJ91U4pNrSESbmRJ0eqv01W66rXq
u8uMF2GOXsgUQAMop2nzdoYWlxEyLl36A6R5hXozmNupmw6nH65vIFxpaggSz2GEFMpd/C9Kift/
FeFSS7nj7dIQ+8znv6sxbMBBHNnaiR0r3oTWxT2xgE+uIaHK9DSQ7EbB5QwACOFXx/tVqnz2UeTw
duvVO5LJkcZ0IbE/RqX2tA2iSAkU6N2HsPyN7ZVfE6yIybqDt/m53ciTie+a3Ug2RBcI/hmOH/+l
qaFxiqp0GT+bT7XASG8jk8oC2lcytAIdWGWDG4eOiF2bfIRUNyI2UIjdF7hBRN2EiVPfaEUQYcpI
GU7sNA5JL0eggCOEBCVJsrGyF9MnNVLTYZB4kn9utLjgkpHIvmFltaIhxIiJ6Wjw1CM3RYe9N9js
Qt22Hc7dubF2YgZmgTY81I60I5Wbh2bcUlocxW61SACQQbLFdpitwhwukCMG20+xuE3FCsMeLBa0
RuSOuoaEiBStAeS8ob1ZlKftzM8e6WTBoDOVBK9bdWoq/FgyCwk0jdM1Y3AbRf5Wdrp7fjNIYuXJ
qAo5hlZ3fSK4ggrr+xgaGXk+2Zb4wJNUJwaGEVuG3gZWZkjLUIaJnhv5Je7xpdkHFUR64TorYKXv
2X6sdIKUEYCa6sq+wnMG3PrimiIv7cVN6dFjS2p/UiNZN8ZV7PZga5/zdP8v0j6qwtksXp8eUuoJ
GltnN/PEDxVdhEhbCTS8UmPvKP6USJMeAuRuFHZJSWudhjjGmSyq3nKCEbBJPfaE4WoVvwcBOXcS
DLQTk1z83HePcKnP8Z8bBPaM3nZdrgycBNnZ0J22w7VTdbjoggMr8HCcpurQ2yxBpTIA/aIJfmBW
kHDujQ52mg783smAYqu3sbQbxht1jgCamwRd6Ql/H+kijYGDBenklhKqPnXa4tzNz7b+aOo7w1ix
oC1lI4FGd+oA0HEZjHp65OyVnBPipC2syJc/0QVJhcknk3ZxctNomzhZgiGZ6OEjLZuKFZf+udGl
qXuUKFTERGFWePwH1Pj4NLCgCY/X8JdoTns92L4/PcsUvTQtDrnqOe2PjSSxFkJD07OmTlMEv70d
kTJgtUpQ9Bkhsfs6PTVvUAsHhn+/ZCEBYiMZJB8aGUGRc4KCEZnF8MgF5ukHSDoLZkVpg84wfJ9B
ZJexKxdsE/dVbCFuizsv5bIwgAxY2hDpaAWMkUq6/xBw4cRfLrdPMUSaq2e+FT2Za43gaDO8yU8H
OhVuyS29XiFysaYhR9OaHOCObHeKgBQR/wbYX8P0ZR+uXGcs1gWr4BkuVxi3COP2iLEO8RSibV7V
l0HUHGqN36IUPo1QYFeGUuTn0TwWvZSNEw6SYax2U8lS3YcPNzxUEPU/3KaZ12psJzpntu/e+h+a
IFMVUQX600vZFQ+ABIbyw7oba1JYMH4x8pLDsPi3VLn99ZwQLmcPd99GXfI3fwknDGKu9xAUdmLR
ba2DsYIwqZWC0Dq6MxnC3xb7CS9+SbbSkHobcFGvBZ3XVmTm2mc/hJEXZQwC9hKLaPcRdC7wwEp3
BfF6C9AUqkPSIXelE6u4OH/r+L3FwErSRe08OtP7koEOTBEmyRS80IdbxjxLnxm3NSnlnF5NRi48
jjoYszjHrNGS79p2s8MTXymD2czteYrNpvz5h599kVG0jKsaNhA7UFk+qPY6nWBrYq0KOgKL6vie
S3exVmKKnw9SSdcFrOKk9vIq2LhUZ4NcHfDm0aVH3F/Wda1rS664f1lN2bGwdbU/1vzxMfuXXzbZ
fbGCO3skglmdJV9XZsAOdlxHy36nlMlMpUBqXw6N3f5g3GlQb4z6zpjd7Qyavh54053PkS6NcVa8
ckzHhsnH3AoPKCS7uK4vSKzPEObjFw5tugRul4t9UyIuKimHsMG+67/RGN6kFrstuj2q7Luauwuq
B8UG97+TKnbKvrAeD0fKIRgJzlxo0KSPguzRPXN3+rhVkYfPi38gCuZa7Bu+oIz2y0yskGP8k99v
11oduN8v8BIrljzgUQapK7KU1Q/L5EicGaSrZYcT9xTWMBh/WyIDJRYgB0JL6bucW5ximjvzVFNg
iG31csOaIcOIDWddjounDpXOJqH1fwGOQe0VIpYWV8qX5CqgJ9gZpjSJ/uGv9ToRoMt2f+JPcdAb
+58pmJpDys6cRKlEEfbD6f2SFQ48nIZKH0bCDirp+8TmDN8/gpRgZh1FFj+xLdtth7A7YzHfXf29
jJ4STAr5WmEtZ3G3oLH3mpuRFWafzypajcK9YyjMevnOWAePlfATs/PZvN+yMqcRIwkH6eqLiaAp
eC55tiC5UCzjtg09Qtav9hQ7p6QN7MmFCsN4Ia3RFdhLWSCVZ4WZb4+dANBp+TfoAv/zkJ3/Q0Bj
O9SZK5s4wWun83QUzcG37dRkkgqFcJq2ziEwh2BJ6DMgtyicTBj7TdDxYyYEwqR2qhiN9nhuBy1D
rMy3Gj/jUzsCRkSmWa5/ktutjhPLYZeKvtAlcYZU7o2wDuMccHodKy4XFvtW9w6hEeaA2yHsXjpY
H8rx8DDDydSftXfo83wn1DHr8P/Zt1mFU+RlFEg3c5gjOMWYpCXNhmZkV9k4ohDd2tQ2sZKhDpYS
I1nNTroXtRrOik9XUeK9YDQ1/Nheemb/6oZnCNBrbYJN2pBl8Mv/0bmrVwRVuHLQDVufhrg+1iCB
X3+l6sSnexpFjgkyL+duCUtpBzbGs5JBRStNfMvTPWuZq7uKcGnPa1Oct6XB6s9NCEcT9iwnezuf
qLo3ySh48dNbJhavvkGwQda1V904lhBXI9GsOyCvPic7tkh5hgm0xaGO/YFHUGOZ91Cc4wXnfcXx
N68Zw96bSAggb/wySw/v/zXKISSLtOsnR1tkVO82z/psjf9Cbqhg0lkjACDIFP0jEb0kgfEQERmg
iPm6lgTKGBSiEMsNEKwzox9/MsrcjFlxH0+OF69ychNF/ikXcyutCdi7WVWHnTOZWEIYE1rZPtyl
MkAwn/03MjUxfiMA05n1O5GcoJX1DewxRVswJHrxZHrGB2+V6N4Q+vaMOuwiYlwuPS+uHDsG8Gqh
yPSNCv3evKVWA2niB4w2ozYkdi5YHa0yQJNrmb/37HJdTmylEPLftrjR3WEsZHKNYh+7ZgKzs8Xm
bljx5/BN+8gQKY76Zn+hlBnUYKQ2Q+3AMueXPWen6yDkie7YBgrpem31nGjxGn9sYWcajl02ddaz
2Ho41S4dAQbhC+tK5WJTwljU81fnEWLIBYG+jYLDMCcnfxLFPmTl967tsNiTs36foFld4P+GIMuF
+3TYBHq3M6d9Vkx8dJJHi+9wgHXx5L8QfutMaw9RqVuFAls8esME62aaJb8ipJoHXEqJ1PGubl6b
RXNrDat7ytMrXMtx77xfuzRXpd8QFqDwzY0gsTSsRwRkrAblBE2uzZ9m9uHOKNI6wpBZoN6AT+LU
0+055Jq3ePShP3UkZCA6DLYSsnkyXqaTzYqoBG2VAPVR5+rkUStAAmh13ULImvPHonzKga2CRx1B
9FCtN1+xEEDoYAOq+Y8HLU3cWlE3NBBzXY00rvHsIaGR6cJwHtrLPYVJyP4/HVqLCyeakWFl5xeJ
xwbVNhYYt3YEBfLe39u41beHfb1cVDNB8ojR4JAi/KufLArDZszFdS27IMZOu+DrOvaENr6IjRsT
fxDt3QnGHjwt80jfCzR7JCGuEwkPLSlX/90rkCllZO1JdXLuDa6BmPck8JplA1xFHdg+3nRz0+8M
Mhn0iJi/FXFAcBAXXGd0d4p7Dtys/rJ51GfcLHlpWaB4PUlHSxoDt02bBOTa+MicP3f0LESA/jQ5
CoGByZ6g+R2sW7W7qlvpxSU+8IhyYFBHno1iO4HJjMreW48Ivja2QjsSs98DZ1MnWY/1AQLjLo/Z
Z285SEZBD4Ilhmdcj5WwkKixcypRd+WPZtwQ45IRHHIhAo2m9apZ9CS1UU49Q8V6NxRyV5Vwn9gA
H+lKQg/foCoa8sIJHsOY3joJ61TwMcZ09P1Ft3NxniVfCNaitIoygQomlo3WWa86wSXdcvOZfnMs
YQqHGpc2hO3NtIznNkfMN16lgid7ZZ27al4oYB2IU/oyj0+lgRu0vFE/wnHzLK89v3c+a2HPbs5V
/nkokryfZp4PRUPe0yj/KiHs8pN7ea6mGPP6b9Fo5iwSRWUx1RXwwH41NWwuBzQurtdI76yKYzyM
pojvP9a3PCbF9mqmmklcJuCZUjdylDSjaKGUPJHcVMmCmwVzVWlnySgnjBQ9cV8wyOz0nR60educ
OtwNTn+hrzOZ3xviO+MCIJB02yir/fJLTUmVFtHytcRikpQ7tvpq+AUDfRQoPGlYDEmVVto/C3Xp
8HnYzufLFcsImXY+BcsLOLPXRSWc0lIdjmmMGJ3U1qwuV01W9QusGbhvfR8On21Zmol51sGYAJe4
ZWhcpP1Nsifb9e4kR3FIIvQ1aUJUEPNGrw81aGoyakXKadj5G6j4Bb2DbOblusDTlGEPV43n2R73
BBwlQ07ct/fiRTLOZkdeEzQHa62RDiTnOpRv8k1lg05Guyzlqonj1zByNBYp3Ro6Y/IXqLmS5PwF
hcgNOFYhg9lugvR7JqGXjt0VhTmURFmNvuljCJwhqn98xW8Zk038wl36JrGFCV4C2rTZIa9/TxgU
Th11HpNGHbXGs4sz4O4y4k+t0/ReB+xEWSeP3MqLNyqf7g9mXP3noX0mj5ih2iBsGVgO9R99Ai/Z
+1TOFhqGksIZDgh9hw2f3uUSapRdhCdiFEpSgQofcxoyvsD+VOmYg0/ryXKEetHTF1iVzvelGnFg
63JIpv/8hPft/VVMh4QRBsQTK2jfla7dEEEEiJDFZQ2x2NSFG5SYe7t9NGqG9mViC8NyEt+Nn9im
jT0wPT+hrwNKRuz/0imjrER0KQy4bFHN6ojwPpG/T5G/wWKsPiHB29Cnqm/7bCCmaRI+z6Q8C2pp
VsXuh7ha9JTp+Gn8tnac3kZmB0hhbRGdH6714AzeNFMz51d1s7lcyvI1GKkP6tPPQ7sBNiLnB+DW
hsmWI6/wgufjQIQKU+/kzatPZ2to7zTk/K7ojksK4uOIOU2K+a2CsOhxhKQM8v+KL5ErA7MbiFCq
KUTyddjKxAQpl/GexT7zY1bEBXLWk63aIVjG1Ff09/KTNmIJr+jCtXbm2aU863Lr4lZ4CuPnRPDh
XNUvf3d9VsYPctcNDXfNzx9r3Nik87WzdycyUXcpFPBWXF5OyfXVln6OhRVyM/CnBOYRxy1E36s0
CurG+8Fls3Y20zXv7xxuuLYXovHkECLkHANRALejqqx06OvguQusM0V6R2EKgHDO4s0C59yZfTsm
vT39ZV7e5KFnPAwedBp0pNhM78O8wwklIMkXR2n9mgXGdoLU0OutvTO4vtiga15+D8vwT8xZcCMQ
3JWgpkzcPJzf1cDDrnTqaFeUc4sW1yAF9SOK71Bw4epwI0oJ4tIAr994hYJ9Zq6m0TyqS8PkokGk
SSMr4wC8bRv1rPsfLQ3tMVKO3WHrTWc+zPCuibE8l1fRnE1DYfNLM9okx0Gu4fXn9AdxpAoM393P
GnFbtU9jhHuOBnwHb80rwBATmuQrTGSKsV6owE6whuFWytlo4Uxe4nn0WipfeCwFISCY0p2DkOAn
a9+TLzobBvIB4jtsmr6JaVAYVEUNpWErGG4vkJhZfzHbo3CJ1RCGW7/8vcsLScY0v9G41yfBarw1
ao0NJ1RS8552MxJfUWF0hTLzg+HyPG/f8ONeSjyKxkMPgdGeiZUz/+5Uqo7t6ksr3SLMFNuY5K4e
fWeQVXdx3oIbeJN6BcHdtKiE39uhCCPaJrv2kRIeY9ivs4hZalv6LydYHKIVm0Hd3GNd7yajwNrJ
MlASC/4oMBClTO2dNiXe+45ecbVosj2FMTq1Om47Gm2ofmNunaoxpAymj5h5ftNGl8RXXK/cI/aL
33wxQE3CKK68qBXqqM3rnj0jzfUSc7wtHx3uAvsSDmAA9i2BorfWOW4+NdJ0pVyEP3zNdS6YTTdW
1ptAqJF5VIqyrqIjnIArMqqos1cSdHJ/vNEZ0XmERpKwdHLO5vff0G5EuqeUT5pTdHfRjmZ8mTAe
E2RHw+fybXTtlN2b0qpwb/ldkxv6S56CuVugchg0IUSwgTG/IqXxHM5cD7+JGHpsCQPPW7eMnR+8
PNXxZAfw48CQLqjLYoVTXKiXoodjvKYy//tN9NijxH0Wixa1+1cnhFXQ1WMgNikGSrgMLi6msiZp
jRa9LL/R7yOrvvytC0nXuTyya4/S9jENN8jnhS8UcleJULe9hSyhsvNuSmdLfd9Xq8TZkACJie+f
o5gRnKXu27pmvJDZsW4jZbwEr7OaHlXRqSabOEZ3qRq/M4lGuEDrExwhFiQz9jqmhgnhApSPUItW
fPUj8oeaxPrFYZGnU71V61WTw/iBUT3qJtSjXRGViv8h9yhoag0jBdHL4jVxqiTcxpe3HtyPup0R
ENcV6h3DuALSA7/C52y59hAdAIsfZkTckvWjjw6cjANGyKlOgOmXLz1NYTDlnU2fiaQ/FLMfdRSl
3C+xnNVyXqQboS1cR5eNGZP+kKqwSHM9w4eEOfJISsDrEbeBsDLhXmX77mthsUHcbz6i+40/g1v6
JBQAQAgTYWbn5ESiuSaM3f0hxOo/K2DC0hTh5xVt8Rt3SMY6n/SgcUzuHFGx4ygztqVjhp87ISpr
q1VFy3Zqqo11ukDQ0PKw9niVVelNGGB69Z6sryLQ6UCTpkGdRpoLnBxWHDnCw4U3xipFlyK/iU+T
6qbaVQEV4UQ0c4keCHC0+NaPDLfb+t2fxpAWhsYTCqX9Jh3jXLNuoPTlU/e4oN9cOsvvZ2n/zz3O
GcZKRNua50eCv4G+D/ODkeW0020YKA4Bi9FMiUKwkO5bR+m9ofo2GhwmYlrklDT3Hnzqzm7LDOWP
NGVMPFzt5u2mRzS+cyYj/TSCSDYZjBSQgd0zoNdoj5IyE6LZ9yz5Tq1shAb+z7k1YlFJc/kLzqWh
9xIMkfZJp8U31LV4QTUHy26h16h8+I2mhdhH0hUMUalFDXQ35g26iHuLArUgGyMhphQUOwqcJ/ft
sIfmazshE/gFfgqVTzOu5m148NEuntAc9b9MhRyw9y+H5SGope6SGQEt2CQk8O++Qn7Itf+c0tfk
tjaRWcx8wuuY3n8k0VOdAd38UaE34lep5bkWxYYmrG4kyxVY0UmwJ+8NlwVm2mwo10NJcJiqm/zq
OFwWnF67Z4+JQYbiU9OT2oVpFFimwsuK1lFm41sfMUoRZpH9mU7QFDe9Qgyq+is+JKD/0Iedw7ps
VFZGEP4j7frnYBsu3hGX/hujlKcxwH/Xw7101fAtIeyVH0JzSWcUXHWEqel36fyhO4YeRTGhabGk
jUL2fT2ZUD/Z9SnUpB3O29MaLtuP8TOik8HDp4QWeURMdNAeiyOz0CnhFpNqdWdb1mu2Bp95HmAs
MzgUSwuPnBar+Z/a6BmGswSE9CbOcWvLHU98UbysRIfIIogs05Hi1k44L9fViS/o8IdnzexuaNSb
FpU1ideMtHpWzFg3B5hZFTz2mxTVmdru0xEmh/DdKAkSmsLPCJxgfFQnNGvDmBkaVYQQUW8lopo3
K6CW+a0I4vq1Ve48LUvwqsyWMNfo6nr/qtTT8qyUo8N1MBwDP6hp1MoYeZu3ehHBg0TrFvG3k9+c
xA4xYMhBlYS1MSZhtdnL7m/eqWRNDfujGW3rvXu6ddmdVaXBO15I6w5yCG5xE/LDu6N0ge3OBlOW
X1U3TKE5EHahtFnyMcNz6YmEUcyOpEHuGAPQCCXhpcKJ17Jc00TrNpiXH/CwGyBVqRaqqs3wJu3k
x3oWHe0ieVXdmfUtNnSo6smX03Y2UR2vMUhmot6sbqx0ypX9uRpbO63uz8sADI7I7MiHmI72WOuM
PbAytoIK6LiQcoD9o8UQNvn44dWOkftsCqJmIGOg3NkjvY9wTPf3rxjb9qN1oxVB7ysXKhh2eoWs
opaS9OsdyIudvCKy/6BGrfArS5mXNjsme9sLpmMf2Um3SXUn3XE+RDhTfK5JOIVgpofwosFEoGyG
FOBXN/yZABmYdhAdZZ8eoSxUv9NyoLaB6uHFf5r8UCaagdXu2wKyQCnsKWvnvDI/GzeVjFpUuz4K
LaBjn3tpF4vsIlR//NRUiHzczekpcYWgBeV9DeSedtb+okB97aYKJvlOBiJZxv7baMMONoyTN4YC
ZjLPzpy79D8Zs1nCuAN1MhosBEGKnX2cXOHuY0AtM0N5dHZw0uD2GJhiAfFihQ8X1k2Cjwz31Dba
1zfyXvqVypB6u65b+fjeoCJmC8Iab8KvURmlG4beD8GOHZc2JOLZMQhpuQ9flgS9UMrfsJmrCp9Z
66BPd614bbM4WNpC9mOMETyOjLHuktS6cYLzJMtvHpeEVkPvPVqLL5t8tVCKfXSlkwNOOVMBHgaj
LdX/VcWJnhtObG/ewnduE2X1GHaOInO8TuP0seYNY1jmdwAXMMC46qOW0fwxdBFcXB4Chp3VIqZp
O2Wj61vOTHqpHPo8DW1EWWHtEn1p482enZtSIe3OFd4u63m3in7q0nUdsJ/GS2SUjIqsykuBhUHP
RTTdyMiXaDseM9r5DCp6SMx83sbuLtL+B1VqGWXx0uWdZvo+oI3ohY7yAP7zp2cRFuENrIn5M8a9
bmmBXYEo9f3DgyNVYgSMlY+m3YKBlBaZ/+KfdoFHEMkCvFzCY2ClDUXEogX2jHftAL6HztgZEn36
wbCXJYYBaMVNHacRD69g7rQd4c6HZ46oIoIVSxNkyTAKkOnyanFfBf1nHuhqzzBDsE9tbqeFoGz7
uO7L/7uj/RtSLBaCDudFWRl4iOQWjnnYQoR/vSwP4NaRkVtOZIF1vKB4YbAu6jiq2tq0pKcAohlx
J+GC4qKC/5KkIPZz4xFC27MlMP0VW9S34yrOzvJ2vxZHOInFDQeiYF5Gkk8di+Bgc1P5ROv1ZQVw
r3wHr1+2ONA5xxwZIdSZhhkVwHCLvGatgbys0OqihasNwNyYfNadqI0Pjxu2jQaH7couZ0Dz5+Dd
nL3d1fHopW+R+JNKzE8EOSaL/KB6kAM8z66zu6kxxtGPNJPJXJzIPKibkMOd8xf5hv2lxJ0UdBk9
TGfqCe2vcnqVG0D5KP5t0Dl/yJ5fUHaqBb9L+Z/fqZugK/GoQddwj+tBKXEWxAcbKF2JBfbSeNql
RlliwWYbv+9bSIbcSwF30re5zvm+nzFfdvWsKDH5ZkhLqlgQ261wbGZW4jFQ0AyPfsvvc0/Y0RZu
SMeHEYBuR4g7Dno894FGTk048B9E5ZXh3ClRXtfs746HML+AFl5PHa4XMTZhtpGLul4Xyq5rY5pE
7YOjGv4phB389In7DsflTOcVRyH3KwiFgBOSPK/kT8wa9Ww8+psDDEr0ro6+5CWnzYodyh4ld7qe
LUoM57adpdfmXCKWN88DSQ6Iqhe51glJOzIWXw89KDrkj27E5oILc6GuIO9HxAk0nIrh0G7QUcYM
TwPcVaG9N327OTm9vtj+3apxuKC6JGJY4lMEDyR+mWuHv92Ksap3iOk8MaDh89MdWGRA1lMANDdv
GcqbpT+J8p6UlzuzABS/aP7BjLbEljD3GGT3nj/smYzP7hBjfPoLOwNd1NAO9frw7/gtbreJTuq+
tUzY1B8BcJUPnxHIi/hX8jjPTI0990zaIbqXUyts/we4GUrK3UV5dDQ8XVz7dlDe+l9Ckg56HPQM
e8n9oV/XQHP0tkz9/z9Z629yvlEj9qLYuvhJVoNtFZlDzL94A+L+5pi9kGkYuwmnJS8Jo90x9yHW
TTk4MTwBo8GIQIGyPopObx38af7SvECsyNgMawLUFyYoV9AGWTo0XDoo3elOkLI2xcTnHWdqcafl
bJjetdmekbGfq+k0j8VgEJLyvplVS3ZzA0NpgiKFZSDQSm0naBKw0nCa1vWzvttzTjAgYSmKQD3r
TOunUFvReGqg4uc7Q3+9Y8+9s8TLPh1soIPqbbn7tTtFtSuAr8Ykgm434Emm9epBgNLRE/Mw+ofK
sC18xvuJ/ZncdS2B2UYYramJ1dVthzPrpyjf9V2hVenUryLpUXB2LBuJAV6yXVk+/zYgkQWdxSzt
5ufy/vZDU1FStyTJfjJzbmPrEwK/KcoesMfs89ojvuqVqjVXQ6Pcnit9qIt4AbYKVsh8j/ABfBQL
UjP8BP5kyhxg9meKD/we4VqOrCPqOffjYfLfEKtV0eaoKQOkXdlm5vc6wOnCCL37yfqEHF08CEN4
MdQ4gRUJt/9sUbFSeUOjdFbC1vCVdJXz4dITOeozpLWzMmfaIobrDn6rr9eXWO+TNWKslOoTvJBb
Pulp8ktafn185RdbiiVnabtLCPTbS3hd8w5F/aCmnDy8JiHowdByzUBTGXTvfnvqV+6fVsUF0mhN
t5vjqVlNYMk0RoQOxRW/Dnuh1CIz4kYi2JldPwp+VhQtKgCEtk9+02y4MAHw3f6GQjI9je7Mq0r7
M62f01OvXw8cLDaNbhXg6/xpS8Li1LLpeTeMS5/EY1LDlzJmeKMr5jltLlkc4roYDCAF9ogO3WuD
D/NRTZDXsLkb2GTAMqTwr7wVsUzFEQyXwybZaCNQdikagIkk/Nnv7zjolVfGD0IDbTu/2uKeUHwT
vtikeoBV+wmTLWk/XCgDmCAhAuhXFfE0M8LJlpf+ghoPcaiDKVxLXwJjvShJ9LO3ebM+Mlq90lol
eXBSwQ5pDRyNHDVdCNscWwI9N0tZdbqRStAjIWfJg4pMLSEGOoQ117Axi9eQBxWI97nvdm2saWne
CJsA5ovsP58eheL7iUw62mHASgyrQdPM0tGq6pFiEydDYWsvhC1Zm63AzMfFhZcb708oK9ez0ojW
EQZrCohe+zOfwjF9k+tAzm3FPidOu7uXkwEDcmMY815q9nyPWLPpcD80heshzelysMwpjeGtp0vU
Uj+vVyEGL2C8v3ZJQ3j1inUEyrUujtbmmaa18xLU5AuawzdMJSpSVITynWShwnUoyAJAurTetVb9
Wx0fN+bOPJvbEWGrzuFsVkaeUlVoIl+P4hi9ND7HdS5c3wljJTRb7sW/e8smk1cVh5tR2Ycf60Yc
qP4Pdl4RAc2ZAdHAue1R12Lr3tGs9fCPbCJjJJw0nUiNsOq3Wc44TXlbA2+5x7FVNCC4kLH+ItIi
Uwu0oZ9jP8OoToBsiGLmgVpKIwOy3qwUx13oCiH1cj7bawG3qCfh9v6rUSfVfo3M+t+eigQrzhvS
dk1LeWvrXDBrJ55ZK5pQ+6IpWAuN/6CE9yAY2UDGc/RrXhie3jr9AuwVAa77oTvuz5+lGBeBPA2s
AqnMNwN9RlJbNlXASqkvtNTG3JwzUOq+aqi0t09rffmdB7Z4vtf/AWgOmu1U/+jPzwIIDN5btRmN
g7Q1Twk8jpxybqxi8JwMjyXB5YQotygUgjsKtiB1XojIyj0slIR1FbZdlep3Q3/VWZz3QqGqdSjh
jPMTW89LMpMNyVBxNrCvydoLI9ueYNz+24LrrA0ILxtjA9nji4BfVlob8pD6B/d2Py5Cn4Su/SR6
8NEpHtmct6qNAB52C4fyGdreFfYVg7FF/yJeNDExoDY8vhOdx5Y9MCMAIxgf07XNmo/qEMdGK9dy
XjTiznAY0ndJAkNM8q8ZWzF4heuB1DNY6lwe83PXS9j5cVgPGdQBvX/2tI9sM2QNiqCdkTrkjyPQ
mTK5krEelH5fvgBPT1lB44XcGZIivcj4OkI+S133mRzccaLSjJ039aYiJ18+2j80tlKl8FYzXagF
V39I6uMZp41Zc56mPukovxQonQPJNSo1Js4AvrQuj8sA3yffwLUxA8XQ1Gmex6oWVNgVMghvB1Jl
DlVFTqju7X1hEf9iUcAMMoXSQR7ixUyWSehIT1nurwn0ByBvAMPC/+tVUBzu/MEUKRVjQKW4ogFV
4jirs7ooyzuJi8WLUr9wRI1nOJivot9rlRlpY8QnfTvjttqCN8bFAScqBvL8CebG6sOFPtfSECpf
uo7hysyy5QnCnkKUrwldCw7dhvqNC9NId/+UWz989NoLBUL0j1eRUtSVIMB0Zc1NBJNBFncxgr0a
u4R7EW7pfmdRK172P7IfpHTi0Yhg4Ad2bVSanvReoyfsnR+3AQ2/vyn0a2OfeQT/wLzzSJyeG9gF
TLSLw6FQyoMkpbrbgYgPid28XMVAgMqutTp13jQdm+n4ePxwR/3dJhEV9Ttl3OaowaCRo6zKDoAR
fWDZmsPSRiDG0vfKb11OadVdWdG+MIfqRqoQGjQ9CWoagR0hF7ajjDJ5yQyWkVNZwIEkzxEEhBXR
OGAlYGtjxRd62OmT5ycHCJuAxPFP4fXPoI2txFdYrL8fChJ+7sbyxMBKQIk7VomRS8IP/FLte+OJ
Txm3d/oVBgEyAQ6exRgFQOrlXCL6cLIb/P6jgX/x8FCVQJ/3Dz8oU2ELJDYF3Dn1yvU4YzuLsqQg
BZTHwNFfYiz1Qgp3jCmh7tZpqHil59QM6vS6ybzDvHCHRbK89xMeNQE9x0a0ixhcOiYk6tLEEOy0
7NizIuMP8fRRDqZ7hkyTEu1Ers1RS6aqTphgeTmzJ03lCdGAjQjGOukXkCiX6nWBnJrh/FAAkmEj
uOOpkK6gaP/sFZxw93xjSYRaiFFFbjlkRo04YWA8WsQ60AfmJVMB2LgbzpfhuZygMyP3nQwYpngz
3kUaap1v75zPSykS2jVzlg3gUahzCMQxm71aClXpfBAL447AuPpK9JYoRTmpE0cwgOP+bSddN4Ab
D4lat3wAwT+wy59haCJJm5243Ed6gybI9wrWvW5EOC+4ZID4IDVA/SCnsPijxknnctixkRcjoerr
84FWRGc0qW0dHoweA4eVRTYZOqtdl6+ZoynPFzULU5VKVLOxv05fqfZ+qqQH382X9ClEyHXnutol
eLdw7Y0kWWYVa53EZcnWYdxnb7gMMLXUPs1PHT9o11EJpd0/WJuqU9M89lo63d/R3gDt0jPReq0+
9s76mBZw1puj/UoK4767NuO1zQV4eMaMy8dqhfLdViy7FwzJCSw7F58RC976a0DGVagkM+mYMNb9
lo0kgxznluwrmYaSDADCYhj2hxnPDGzryfo0JqLBD5XqO4RsaA9Z7Un2RLcApbKaXMSQfEJnSpJY
u500vlt6ZbgMkUNiGMJyQYAaltWVMhYw9ubwqn3hHZ7orrPZ7lvgNcEt59gp9C0UayRTGoXedsu2
Fh06WJS1raEPifmhyNAy/BIm0RJwzgiu+it6YLjlzKxMFlnCMQLWkmePABT4841X7v5PMDYCIliR
wCXp3QtjwWJhFAQvaOxvrtIY69Et6S1o67HKgRSfcX3RrhGVpnvGP75YsrSCYf8hjBOcsWPa9sja
MrO6kSFxjJ0BP5vPobrOP3mRjzM2TzaHAUTstkO/k60NuxFwcj+lBePPT0J+0ZuXVIlD8NXYIrT0
ySjRHiz7oTw9gFlE4tz1dcuJXRZpaQoyiusVrKkuj72HzfRSzZV+ZGU4V+4zHwz2Evert0WCJzuo
MAj/xet3Ddr9lPIFbUiDb7EwIjwHZibSsuxsdQ6XWcCTcfo6CT4Ku7pLaT4496VZtf5FiFbnn68l
Lb/iVC7j3rctJqWbDMAbpM3m2Fd7s2LxSbiyR6H3fmBJqlYB8ZVzSSPM9XDqrprl0stxgx7Nua5z
hnjlx7Caw35LmE+Y873qbYQJfRhAPV2R8pZBp+MFZub6DQkEVTwms1IrNK1a5lpMvGL2LkOt0OHH
pbvxjjhK+IMF7EIFsj+na+BJ1QwqXIejWtprdVjp6GlM0y+hy2JIiw8a5OVjMlJW9y1c2w/DxbA5
plAXu5RUW3vznPzEv1555Lj3+ZCCLZ+vhJqC6t0unDPW2K1M0uQ+ra6XXWQ1qwT4Ep5Qgpa0/UKh
eWG4CDKvDguHxLbhc+0NPt2m5ycbl0Vhseh+GrUJALcufN029zptYnjQsXcn3N/Kr5fTaixV+DO3
smQi0/kXJvCUm000kPLqUqaD8N5tNfCk8hIsLAGPPr1UGcb5/FsK6KwgikjtWoiaM0oS0w16BmZX
eapCWLKgditUCV4m8eyUyLlUPL6eijKvnOgHsofO0Pdrq50XtYTbJcVv42A2xZKOpDu3aHiRi2wc
kj4k4Iux5jt4+wzuzHE2LCpB2C4IGjHSnbqo195KMehZw6J6zsShjUIXd853ypu0+Jdn8amwmkhN
6A2JOlL4MUEGwV6f1dC+NDzW+kdWF3k0lALnUF7Yn4w1Yi56qwN8iGIk8csK068CbKgYMyDoJ6wY
lqd7VbMcKqdQGavz2t21CaB7IrfBLOCH/gqTiRET+ysKqdR3oNXc0Ek3qkAl6Aet5tgUdx2oQ57A
of48uiMEmb0SjZbSPZBug+K7dEFdcaHcsHWEyzqDk2hMyog5uXPDoNMo40wmE6/3wFV/XYz5Nvcq
NV8iVhCO2h1TrFEHnFxTqzSNMbGfxvh6RWFAMG3sz3SN8DO8IfbDH1KCRyyMBx1XDDN9Ghn7u+6T
LfDATVcJAVQyKzJ+BgMTWswcmR6qC3ZvcLXDS8bmYGezs2AgJNVDWCDU5ZLNArQbuZNFQAMYS9zy
oW/7OKb62xdGgspL/dHWwZrZcvC7t1Rk7K9qyaslu2rWpX84hD0S5SYNvgElcpdmDbfsQBN4d7Vd
4WtI2qsO0ZMICz6rVWP+h6dFtrLXCCpFQ7nvNdfGAxPFUU0Xaf7tX3RymZCH9jB4y8ZLHODWZDWt
/60JldNHBbpb9IsN27J1Ddksm1ZK/SzSnNWdD2dOZkWqzaMnk2i87UavZMEOztre35evq+HqWhMS
cii1WwsQazqH74eYwDPveGPP4yFNqzP6WkKFDoU5w9nZnyz/sbf8vR8ZBD8YTPiuoH5iDD65vXOL
wzrsqAoynhA0IySMpcfrEDf9h4RYBZoA8DAJVHWu7GZjR0gAIKbNafY4E8ymjcERpkhfXnO27KRa
1kr43IG6viZ86OZqyylg2n9YzSKDjmgm+3W5L6WWnH3kwQ5l2mxe8AR1oI2qEaWttbSCgwEvopJo
5MBKEsrGBYJwnNFS7rPogoUmD/CKdZSi6uha1XoEF/PVKp0dRQB18XVl4DyTb+TRTcw3ojbCmuFz
wOVeb+ndZflQCVX6VKYM1TIedhH/1Advuv4cPNwY2K5DC8w9/RNuHdycelguKrLnpSwft+Lj2Vgr
vF3fLmj7CnqKfsTeUNXXfFH/pANjP90zZDPM++L4KGF5WTtiG67r3QAp3/Mvr8TBIWHY+WI70n1m
pflaHaYyZVq3672PK4V/61uFt2psEIOv+Vhum35+rNNqHOMsugNbj1kzEWerq3FuCafhojKpVMLP
oYNXJ70+UFLydLMPvESI7OHl2MipbOrTJVTmSJQgk699pPb1R2siDRKSMPNtwbIkUyBgLQaKKAVB
caVsLPPvoTIgyc4T0KYSLpPn6WiJTCeDdDQkAhpQyier2lxTYbzcuhE2jB+upZmpcApp5h9JEEEK
r24ziPrih6V5mpPIbl5VFCWGtgoNqTav84sgTRSscgqSaVoiPrviaYDLwarZ0+A5Ez9+3FjR8bhB
kcbyDOQ0Cq2wInYFsVbOB8yLiwIPcEmlQ4eivBRfNxA7LsraPPcYJUrbwo+Po5g24LKXWEdjlQUR
wspJBXJ6HTab0lHTs8M3TxGpkqZynZT920jUue+SUtUpQlLoBoDfsk3goT4Jla1x3MGTW5ZoBFoX
KbvoqmK2Gs1JhLBKe9GEmvWFGBn0M5TWbMNicmq8sekhx3Ntb7gNfZYUu9UYoXNKAnKg9s3lg0YK
36nUNS1Uz7Pv0VtBHeYO51FNkicSiiVpBjbD/HijBexNTWgw/4sgSzH537FmT+njU6Ivuw4fkJFd
Kv0NzcTtLXnrfYMGS8eqtc1aDyfhvEBqaA2zpepZVbDXtfFuuLxlnfu1OYvg7r/V/ougeyCKwNTF
oLX55VowOxVV5oOdwcR/pjl5Rb/Ap3qw0gh4Gu6NJFniLNJueND/Gw+aU8WbtYwL7rAY2/EzHNvl
mHCE+Wkx2JTuZ/CKlpWVQqz4HYbJ1PLgbBaEQQoMN70U2MU6Nh6mQ47zsEhpHnzd7186V1etPUQm
h3SgAOuMYqhg97ZNQ7bug7NjLnq9Ct2WEvCxbStFhqx8mWWLW02rsQt8AKTg25cmmnR6CNCnUyTF
VgH3lpTxUlU6fZJSc2DKhcoGyo3eq7Ty9asSOeri4F4hJ6qGEpV15SslKRWnOOYxKEvjjQiYqfw5
bIVepXm/mKOlxoCC5fZCPrnpntL5DLeUe6C3Ob8nIDJIsUm5ur1lNwb4edmamuJaTZp9STyA9SCD
X85/HjfTFsI8ShVMoYd9JnyCnVjfnmNsDsKsDOpZjYb5kHlFIZRISi0+Eqb0AjoC0q03UWAxEAOV
IedJT6DNH0b1+r48+wgkYtRwgZmec5JPVip+b4eg8N4jVmpiEMp/fdAeNb97hM7meb1v8nG4ou0t
wzz/MSB/DQNbL9aSIQCkEn8/OpcnLIcyIrGKWvSPS3If2orK9UrlhsJ+kTWc7/RZ6nkhAcKacRAJ
F+CnBjYW7OmnrGXQ6nBGqtYverNfvUmuOTi+J0Ktt4s7WLROhNJEEedVfAJgiGnYEyjMODfiTUz+
/dMDML6UGW4nB5yTbHQUYEY0lQJ57M0+SYid4m9YHEgx4fAVlaxpIGuVNZrEF6ibQjK0gPlfLIbp
mp0+EunLQWsPtqyKRSarNJE0/fu9ENswq2GJQ1UiixXsGCw+6pYNzuwbtGCEfRJMUiJ4NyCS4dl2
o454gBDJngO2CO6uFmkH3YU7ZfMZsq5otZciQNATEog8FgnpDwYj7/vCXBJ3SNm4LBOo74AgrCnD
QDDZrGzkXy0gVMmorWTi8kZytYXZ0bTgkRfqZOGPxe4D6X4tUKTEHR0+jxQxi77W5zHrZOysZplM
FlBstxxnh/ah2aDtv0JZz07p++ZR8RboffTmzu8my+3CPxzgekt8vTILLxgC0/NgEEtLp7CwaMDZ
khMltnyZ3dL4pplawL2XZHCISLIVTFVURlyMywDeNDJ9esMNrwT3jKCC/c+V7KWZlZM43Ee5yEo5
OxjC/OW0aHmRSladGF8nM1bl1NVp44QP/iaWBWXoht056gtdT1EpxQzpZJRWnyi3O3LNUjp80wga
V3ZgHldBLQsyX8I4wzT8SL3sU7kGziyLGNqVhEDsTfusvh3/fbd3vxyPC1JjG2HY25LyhoZU5Q2A
jDmXaO1il7OrpSqKy8MEiJ9FWx0ZSyJ53vcOwxvrlPYI/CfQ20sqbAbZ5aF4+Nb/6B7Qp3+vy03C
wN77fw4BQHZJAF9s8fdxWNvD8V1s+7U6eun1xBErlM6u3V2r3CHps0x1C74bNQu/2/U2MuesavQn
Z2EFBPTb5h5q/j+VroiEVXLKd7/rfFHjRJgtdTMpCY32bx0lC0LKZ4Nu5eu4hLygzRPfk+VyaS7d
vCJO0HxGnmxkMtw1Ux7V+1xoM5M4TVLdT4C4Ts0KI4z5g+/6UsoFKh6zkEueRGD+8/5nX3LXFa7j
yNzU/nHmPtLptfTS1Q5oTCNsQUKudMtu+StwaKlq8QxS8gB+H+D6DNF4UGuAzxewn62zciXXED30
eMkgR8hOccnuxOFf22Ujq7jrb4F1i2uaq+PLApYY883AFnts3Z80iq8M9zXsl7PuQXeqgoqPwfeV
EOSGQnRndvriu/oyPuA+W3mqS0/6AfoApmtHuF3JdmoiFx3ZQvRPRBqsvDrXB85Yq4NFMDNIg6fb
/aMQSBByYtEy0e0kCrrTCGBdRpdmoaO6B+um68mQnI48Bcunpk/sT1LIyEJkbOeh89Ea3+dTCdbn
PUGlQDmDHPG/5QEjOwFxcwsWsbGw3ENt8IxTJmy5J+Xx9yjMmDNqokf/rp7/MTWy3tvPp9clUUm/
hqzgO6ziqFTgqdNRRyRgvdssXFQ0MRgX1ny7NCT0GwCKqxTPpLarIlazYkZhcEUo7ihN7lvKIufb
UjZ7NWV7AkD4Rh5ekQ3/rlImZ5/l2XWr0OaqShOTn6928LTyJQxvXDBNww/Dls6hmbVTBgeDAIsa
+Tn3WiW87hqpQ0Ql95+1uQqiT2FXjaby4PAv1hrkXIIOm5emOteVU35NP545a6F5Bpv/uPwFMPwX
F7mlNLE8viN5WOmI3DhPCFyeoSCmOID6ElsnlNtmvRWf9F9jbYPk/LY1zI9RtZs0cOEQRKYUAPBG
1YTV2mnllZ6afJ9RPsqEDf06SMuScs2heqEJNClR9NhIExIBYdjQeKarklgDzWOYwNLImA9y4dlu
sJYoe+i+5/MhxyR/Kvtb6TxCvZByueTjJChDp1C5qf7dK91C2EszBthSxYsg2AV1EmXmRUcH1eAB
PWXatOwVEFbvnYIpZuN/8SrN3fXn8MmFnAY+CpEYpt4XG6aaijju89+wl7O5DYC70LzKnNxxEJ+z
+4z2/DT8CrZP+3O848mkB3FdclE45XFKkw4ubhhqYWSrOSW+MqtycS3PcRZqMgQBQlzp6VTTQETG
Y3PKGBLklKNDHe9QUAlBsFh8/eK5JgbB1obB88tpXZmT+X2dDvrrK2wrHDZZYK9zrbL5wJu8YAXD
cE3aoke1ln1YftmJabNfbNCaKLV8Oqd2s+u6qJp8IG46Bwc53ZweIGlZ1caebCY/evQ8YYqdkq5R
NZ+Wn3eYcroUlhqKBuTvii+HS1mbljlNzvP5BvBap1wWlI2q4/SuiOkc5ae2sfy7XLBwVWgJcfTC
V+L8v/YxMBKw0WsLzfIQDJ5LslslJETuuK3ER2VFV3Su5Pd0B5/QMRgekzv9NtZOuIkK7WMCfHFd
1pGhZJV8nj7UnUr+xQbqrke6RunXOvL8aR1AqK6v6C3aOh0PtEXlVng/kEQ6fW6HTzzeRYg5p1Xd
VZlc45JOo9MUjy3o3t6zxQLrOQ8grg04kuO28QkahvI4SDBuJ8lN/FjSPHr+luECkishQT/VjSKu
8rsF8UVVJRfZkUk7b1s9MnRY6i1F6c4VMdX8kgnSnHXoNzM8wts5GBjWpzR6NCOTuBAiNUCJWO0N
Szbc+lp2a7v80C6BK/jkaVqEO76/xfyIb5fCHykg2I8tA3ruT+k8FQ3w09PBhG/KGtnQBpS+/5Ig
T/KEPXD03/9P8sgBKzQnQexIPQFMHADZQwaCiwL5z5CGloumFgLZU94NNWmYg54hMHltukAwHwNU
7N0bR2J6ByeLeAU3t1kY8/5TlvSKarK3v4YkTI0eFK1g/VTuWl9FfY1Rxudns1n5dHjyNUvel/x0
QcHXL8uAXUZ0VKrMMvDZhSnF77PNuQ42r6JEW261AArGbSzw++ZIMq/qjBA2db2vnyo3ot/smYpT
tJlmA3mkf27Ov5z3wK6Wkc9OYMdn52mko6s68IZpAwG6liRIIX1chXUDPOA+DVLcMWPKseS0sioc
OjhcyroDDtI2vBt1OKEtaYczohdORAG0J3ri7G7izjJDKNjKABAmf1Wl0V5AebiaUzq9vfJw9L90
HFePqxivVuAJScH8Y+dMJ3sWT5k71RgsNnzj0QEoDjB56A2G3V5YKOIuYJ1Fghgumw4M2t/dXmzi
FCLdpEdqMdh4vuHu4TXN2i/4Wkm7Ib512J1yYIcz3y6YFw48sQgRbgy5aYR0nT0w5PJoCEQ9jC74
zoVoPXcGwgPNryFwbIJOtKSeb3ACKjDKx+Mwj97zXJ/dM0iuXDJFr/BTqxesWJAKX0UzloR15oL+
uXdH53ydqSxaB0CxuVskO3HskQlvCfKIivIJWNZgids5WMYJMP15Dz0rxIkUv3cRCuyEu2jn6n0K
bk4imotD8HeO4U77MJw0tieltocz0UdTgHMtLl1Klk0u+MfPYYCjki8j9sOV7MhgJso3Z1olPIUW
MLimBuPnEYycnyvigcbrMApDS+Z3wNQnQldR4rdFv4a73DAfTzGKqgn5o7AyOEknaiDXTTYRZzpH
8pFvbpbBTndSqCUIJGXi5BLZpKeYZMkaJFYd37ZBNU5HjqTE6uuYoyJ2dI3JJhC476ebsabQmok3
vY0RXkUn8kJxVMkI9nSuEYxn+tY2Bgx5qSMzVof4HtlLLGDlLxCzb6mLb4CIMbG/w30niUMdvzge
CVfMbvpKoOfURYOkx86cl7WC7wm9hvWwluhfo6rzKCv/5KvVidpA7ed+K6aA+OGUz4CzAEpo8DR3
7hhbndoGNvob1AdIplVoKgXPjMUYBVRvbZZWfWIbH7d03JQOYJuvSpYR6iW+U3uiVzVcHqVZWIEg
bcfNtGew3+rnWg+fSgwd7jD8y/A+SpuyjwxKzXWpzWVJPrNPUYeE5zlom7VcP3V2rBwhbr7PY8zk
KiUYN7T4TzcApBNMp3VLZ0FCyTdLEtvV1z/oQM5aYy1La5qqj3hmsSCoowCgNuI/MdqO3mqhzHZJ
eq7oQphtasqeY+HcOsmpgyq+a3AzPVcIcw0vIkDvFFYRsJkHIwR7pCbmbYiwO388chOzNO+56h0P
8bi32yM/p/0J+Q12yqBA+DQPHNOtuLfO5QjKozrgAwOQWcg5L85HbWQezu9Gn7A6GDWEgFpLmn55
Xv23o9G6c75GI5U+6jBJj3z2OZ38djJYUFOCyPIdxA31PaVdhBN5adoWi+ETBVeG5JacZ4PzwUXt
bjCod3fD4/NSoZSDaIwaCkprGepfg3hEasQXueSrX2d1edcOIZBg4PWcNXxQV1bnF2KNEj3cN1cj
KEKgckfR7bhHL29svVM0nEdUWD0f4OOpQDhlE9ifvdFrjJkvpYeVpXplnALsDNMV3o+c38bQ9sd2
JttNsaLZ5TUPc6QYTbgofyVNCRRHt9wncYne4MqTmSO285MYQoYKHFkAdB0jK9iyyXvbuGQklOI4
EwqZYzFwlU53J4iEhYyk6l5STw/s1nZkrc4OxU33usQnDP53FqcyUpbIcQ+TAeeaFNIfg9nQ5WYF
p8nx8LXMp4crVObjnf/iHXfpolRm/GtfUWGxMj9o3BoksGpiKRODAjZ0nksFFMRWO3y3+Z9EyUHg
fC+g+48F8ihglEPcm7lUiylQ1JEqzSfZZG6vhf62yW+4z0ertmsAAS2rhBAjJIWcTskcON+VotEE
DoDODaZ+oDyIN2UQFsVIfMMN6zcbArG5nVIbLmg2NxgbF8H7PX3afVkhFm/Ltbdq8PRthN28zQZX
2Cfqmm1D9lZwszzV8ne464qq0Xb3ZDhcR3BIcU88QobcjS61icgCe/+JQwn0EplOq8qmWmOdR+Ma
NKvvkvZm859ahlfVhsaE9mpqMnDUmpIzLecpHPHcnHzxSlbDqLqq39tS5liOiaWEiORE1I92wmmI
ebqvSq27BXRyXv+6E7HfOHRqj+rStmxGG56WOV4ztreNxoGU6vAh2rcgA9uGAch9wOUkXHI+BIzk
Cn9pG+DqRVit1/CrLKkDwQdzg63vdc80w1cSNJZFQb3Vu690EV+G1kMrpFiFoPPJQmfltHmAdJzq
pWRr4rj47L1L2X5KCJeXpL7P4RhM7Bml9+pPTXL/kYuoL+9doU5PzPDZC+ErNf4l0YWCnwzKo7fu
Q5KAd4+4FH9yhiNdSqNvoMckFVj9ReCxW5fySITiKSQrXG06fpvmdybKN+W4VZqljL/UuKu7l/Li
zvz/hdtwXEpMVyZa/4MHBVV7niUKra0dfw7jJ1gQLJcg0J55SAIgiDeoQnmZMzRer6RCzfsTthi/
P7P5QPucZMik8iOk129IdJh0WSz5b0VRQoh+IgRZatWvBhG9driIi9Umu0MNlwLos1cS4yUnM33t
2Q41MYlwCPGkeSVDIviQvv8rjt0dyYAulX8oUGkZLCoFiDAinqqwc2SuBcqqhh5QGV4+Ka1vDDVu
WfrM7+4QzvqTcaRWaroKJyCyCdVha9AKrAH6uCe/TLeVzxBlY+rvonBqkhBCNksPaebj+ZxN39Ec
ypO1OXc24cXZZlGFruwnSaXts+2RyfckIt/949G0WXZQgO3D+rk/7Xfo7alD1sCEN1dcIDaFbYwz
Z+n64Z1Ggh3CBxbcpwQ/p1BJX/QGTEgCgv/AwJU2sWdbmM413toJvNKuAwRdt3ugPKlkpZhKOZKD
hYNGnQJdhusbqZnHZhKJW255nLOnf5V7m/TWSDQMY4KNw5c+mAeE1Hdi+oFZwM0eAZOlG2RGOJnC
Sxg9Hbgfo9G7Hsj4cu2is1wLGqwSIgbXnDLct8XAjHRHOEJFRwkiYtT6DMSdYPzW88q0v3lxRw89
UeV30xoi2IGpTVTBaHadTSrKVfog0PJaMiGbQoqyVwlq47nG0al5uxgze3VHAWalfLSfP88aGaXE
PZfmiUVjpN8on4anxR1x03VnfF+Ivj3Wlx1jD/SSEjl9212wRLORXgCJ9DPWT6eqoTX3z0O/0Bs3
qNkvS64OSBphAde7fM9HIAIpD7UhMgzkSweM36GITfOAbUbagYyikUgww4ZXd3yoeSXlbiggDOZQ
lvCQ01Y06tu2wmxxtKtHhK721men7aRW04Mkw4mxYOwbgLA58HE5b6vP02o7mOC/4IWqf8qDXtYd
qRhNwfyt5A62v6IpMs3Uu7XcLXiKdbdJT/jwocKemnYXVOX6V0F/dJ7mTcBiddT+DZQV5saJLAgo
S5TImGJ/O5yvEZOP99R0PXOOz74Dis0ULh4vJ7CiwstRZrweFOryXM/0c4H/dlMElRGKsBcRoQuO
c6Q/Mk3a99ryeI2HZGzY8PT4XAB0yhnyvtlXzsp/ly+Hm7D/xEQgw3sspB+xQybB6FEBjsp1AWBv
4JS4WgEchUmgdKowDYCC82wxsmiJ7GGCNsy7urMnq3P9fIPz0+Ggg272Z+N0GzK/qncG+nTikiyu
yl40jlWaVsqsps/jWfnk5M24fztjUhMRwjMvZYmdRhfYKmiG2cVtXvQHKnlf+XQyxc1tKifdKSDk
deSK/FqxPlRSgxCRtCW5Pn3c5gg9hd2/mKAtTYauxsOiCWQ+sOfNC+jcGu39lGpGGJaOGirESckt
6RbDZJHsq6Lt1ixQy6Hv/heB1Rurko0t0OoxUNKAqr8fv8XmKF/pgvi7Gx2QJHP+mW4m8+Jq4hYX
83AweneGBv4cDXnyzBvPKxEvzSzIxZB05gak0TgZhjCgu062L0AOm93XNGMftCcgSNv4nInZEF0N
aworUXuR3Yfb3SPiSVUpvgwtbV4oXwwWvHBiu89eN6Ie/+2fKF9wYY+V4IrUhaW8CtCstmcFsVha
+WzOsX1ih7iC1i/aFlgPOKSpRsSCLVLl8ax+QrOn+YYl/4FKi8jcklrbLvZPuBmBwLY0BkqG2DZd
Jwa/wfyVFCQE/Ay3Yf53DcFBHU+6XdpkpR7gwR3tOB8fyZohQwKeOcNgAQ8Z+5eStSmobYpGVMzH
QqSx8TW97TvDEKHmAVdxZoyhHZuayDalXiy6tf8cWmyz+nF9Y5m92AyHtZljZOeBR3Ec9aLVh1h9
+5pwhLmyBAhi0MgX/IcZTMIMTG/H+lx6MLONPcF1+qbfR3bV04B0t9H+gpbut03K9wA4tFqZOBJm
kw8pslb7qc2wKHSkMhkDHp4w+2d8PmKqg3EGgrdxGg7og5JL45tDKyBrZmiagL/XIW6Z6R6vMtME
QhAoCPGg13BPCn6EY1lQI66rHct9WWCZ3b+96cqQ8mHdJAm8mkO8Xf9QPBJ+8joqqrTMFa129zTM
ihuRLSQ3bRJBfbBxgl390pY/RnIhW0Wfw3llYYWmWe41rX6ucyFOa4LXZTfXdXU7TSv7gyHq/QzG
UOGMnmgTF3eLdaGNpCR5R4iw5qeYAFViHisW5XYpEUQDLcqyyr2ihHvYsZAbW32NL9iulcH8wuBP
wADgXN7/Hu9MJmHvtQZzTaoaM7EzsbgPXQPsrARJHTyTFzFbodZOG6NWecXcJYjGihSOdINwTDdE
g3Rt8ZxncpGts8sHTgYNpy/sAUb2BmCuq0BakU0GMSM1FxwADUrVtjEfMBC7bfE4hCUPS1pSbG2J
Zyy0jmaFsEY8KkQObUdASm6kw03wgAhAbuFW6Nzrsv1wLOSNhCo5GomU1OVF1eYXA5B/kdZ56ghP
UvLL5v5dH1lbkWR6ekMfJwgDF9clwH8FK6ExLyv63PUgaG8LzdRq+pyuks5bfyHqQXh5+Z4UL+cG
DLID42OvTsBJs+53mfVtQM+oRnZ51iV799yru2wS98gvZB5ZJvm01QzGIx+9NCUEV1e/Qpr7GyHy
xw5QaQEyFoQwMBoKOev1NDru9ns2e8TJeCZCOC9kGSCcgMYp64nMSiqu9FjZ64ze1yvIAg6WLeBl
Sl4+sZA0dj4ytFaUakBsWMYt7wrTk8MQHBLU03SyitegDgVB0YyNb5EEtmEma97saT2sqfo1snql
4x4yUPU8rc4+blC7jSk4KcTMDBXjrJmwAO25E+4Z2qRUY0JPmcA2X3LaETI1+wV5jaccyzMvs2rz
WSmcPZnH37+TWC8dNcvo8gSGigCMrodu2ExnIrJ385nNjNN8k0Fg5VGihYCQ5zoBOkvvdF/UBszd
ZPyE055Lmxh11dK/RTeUGGMWMiMzGCAzCSSgo9k5sEezWr9GB3WV0TdAhA1ZHvf1iGH69i1sdVn+
g4S26NM4/qz1yozVjYGbXzA1YyWRtldrWuZkBD8bsZFCcewOXLfLnZML10/uJ+Hc867TKUX+67zD
7QsOC+9pggEzcon8QWa0iNT+tsgDvq+dPnyiAcVSKpA16+UlWvn6TJn1+BZZ9bMwC1X7a0Y3iAhL
gwu4civ/70caA4exuZqWwucXiJA622+XDs7MDTcBlxqx8oJqttR3OFk1eXdsy7iRWqlEuxXc3FWq
xMVpn6Pg9nQwhFlYp+dkyyJ+iU1/Kep/gQlowBkGnzqPk3x8q7PSWAKodv83l0n9tpmVS0GIBGEa
6Wq5vM2IzrngR5WcbXg5kOtXNjrI/dE4kU/f4BwzRbqQwgTaPKW+eDAR5y/XThdvEavP41LmbS8g
xjIDUnjqXfH7QhXoaQp4bKjDHHt8gwrK+w5HEW3Ap1KNhVLZjdldE0sHanzmRLRhXoxp8uCntfLx
2kqfghE3GSkNv1fI46sncdDY59dblrbXqaqhSIMB2ToNGx7RvguFql6tGLXoYtsyLaH7X3S7WEcH
HvLoY9tQcRol2IQjjlNE3P8e0H9iFvGgPbgcjWnIlXZqvtGyLa6pp6r8mgHGwP6ICe8RQ9DU+dZ6
F+irr+fRFYDrU4mi3BgP1gK054OzMAps90kFRFEFXylsY3qJLQHoE7WVr/mH4+0maqM7PMKSvbCh
9HyCZUWSKzyg/cQjofqhbVuZXQxEUWLlROHprk44F2qRHb2iesdx4JQeVG7Zv73sSYy1jBB+Z8wQ
Ezj8H2ymJgVO9jPLY1hNVPLcsPNW9zSHglv4G8zVxRDqu08VvCqAG8frGGb4fzmedfuVluMNT1PB
gOs5i61KqtBKtNveR9Ogt64W70SoJfXxHr/aWD+k/0uqe4dQt8vzv2vogO+Pr8jCiTENfDUCjhkD
EEpxgVBf8gaJ8yCiKeFvamo4n/fCzB4w0QrVHYTz9zXbaIPtp4//OEDRPFX81Hz5Hs8sksP+PnG2
U9DF0FRNNj+RXSxfCTT3Uk+imbhJpW9rqeFlsZmk6//KxjfDOXJKBg35I4FmSmZKlmOZAH4zTSUY
x6CCGljsoeTX37O67gDko6VRZwyf+z4BKCJOtBy2mdJ9qT11OvJBiIMMw0++WtCQbmMhxBk37YG9
ePvRLDF/nbg+8HBDlS+ieaxnBkaUDK1DMJ3pXN92btPBl4+SDwm63vvthenFYFnCXLUB3g3k8/4k
nEi68XF4oAmhdQ+tfAN3PAPo6rV87wFDGsKBHxGU90xnYlxlrpryLVWqa3kzaXhdqXDHr6Yd7bu5
GvsApWVS3gyiV/2akULG+d+yus2OKo+w5PJOBnCTvPzvv5PTLvlgik1ENa5+YYxFbTZFdF+3ujgO
5QFnu54QmfKvsf50EZrUb77BQfB/2BiCpOnph4knJ3voW/nVDrKCWpY9GD9uMtBj/uT6oiUT6sys
6F2NPYtrBOA+WOqCXVNraNJIsXH3H3W0TNs50A0GWI3NqKfHs+VsQqHmldJPXQLaxCxQ5inYSXbk
mf1Vt5lVqRYaYJC/Bx3GgzJLtONIW1kCanmOGTQ9bEc6jrlISt4OyjjhBC9Hml+3AgB/zyCJxdlL
T1QeQu8puWtN9ClAxqRb/FsKEHrgvdZ9g6pSpdf4QRInTLFXxqRJsbfAYEJLxd3zN/2JAXujkyOc
a8NJVL+WIO1CY7AXBom14BqG8qTnegVExFJkX5M+b5KDDPttl2wwWoJvBl7Atqo1Bbj2xkh8AtGi
ulalXE93m5e3V0QHGyKjYw+xlCxW9uQEEOubc/t22Hz19Cr97jX3vvp54ZdSKMfxDJWDyNNuTMVY
OAflX0sZXXnjUSIqUQMuiYdduAIRwNV7viuuZEfPxCvxwNMPXRGAtCgHqBvP8SHJ83jcQMzsHv1k
cdvnfRXPzJdP9AiZH/FeH8bruFbsuihrPyvpjiAqEMxZOhtNTXxrxhsRlNNN1E0OsTgS3kPQWTgv
Rkw099HI3gWT5WzmVPIudiAwQHA9fRtQMMlR9Um5DOzWsO6BDPGYmC4qfxeYbiF4R8vb4nO2jRqL
9SU/z28A8vaXEqJBKVh4+4tS2FcRFB3LAadlxzRGuM3r/aFSQ3Q2FCzmihHrIRhNs1sAd/nKzIXC
44m1ZbyuRmAatFrxfH81t5IXypjAmJnrBnz18uuR/j34usdSkjC7M3EYAKkZb6mu5sQy007/eKH9
ZPWp+LIF15I+76tg8N110BofbYBpZM7Gh3KJsGMS0nB6IfYyjMCVUVfD8cf8zhaHygDx+M8hrsga
JAaJbCSFtCuSX2nJYWV8yKt1XMHstgCUhtapdR6L/64wJVVaVKEiUNl4+zaPI5r9bVVtzs1vYVxF
jFZJpyGlx0I7XhJ6In5ug3+nSmGXUCc03rnRxY9ZHBJSXRIHL9ZM7RmUimOEcSB4AUXngjJhOdkl
vWpiCQC6WuxOPAYq2AqzciCEPtGp3BtTd0Ii3R1BwyKyCJg+U8C/FeJD7Uve3M61xptVEEfqeSRD
yPE/giMWwf6uGPnlYRL0BnYjCrUPRFW6+oKHsDX0QvI311oVbeiowlJ6gccfeF79VBP1V+/uCNY1
4T0nQJcnxFVVlAGq73/n7dk3dL9Q5tIV/WviT+AaiscCMZaKpG7Y2K7EaCrvBpkFdnSsKrIBekR7
QNzza7rsy1JrNxSuAMNxc5MGPo83TvOwXlOvFZggwRIwinD/fvWz9mifUVdTaafej1hDsx1kYZZ1
l1vbiiZP1ie2LR3xaaUCvvShXwdatLWGRoLKBkdBU3iwl0KwT19uDBxmHsKXotXHm5ylpCJeQkAi
3M+4a865Z77RkaVN/MrSQbNRM86i4glv8hh8gfrvtVoV3gbRavC/QPSp0/uJ3akgVBWJbTSRCxkl
iPoH3J/kOulQUJcklwj3hwQNdzaBM9hreAxw+pFd5+YdDJqJ4WEVfEso/VfJytFmpamvNgVCZYL2
ta4l+cJ5MIvRg1xqE5Ldk8d0yFaXM6da5KHxvA+p6jbq/c3sEElfq3r9Rrlw06E4hI0ObDvZ9+6t
ipBIx2B90QECtfaVRlpFYKUNcUE4Fm6+vdZKMEcCdgTbiiz0LKbsq9Bu0Hjo7deZjjX34r1I4SsM
8ej7zUpaVR8Sc1WirxgyP4zCR8Lm6VCGTD1zAVkBeD3xLBa/48Jzct30w9xO9MSuftISK66l9O7Y
+ZCVsXivZ0VdKrPMq1ePRkz4707YShOtV7iZpppz9Z06Fb54qF5DYcYGoT0/2bRKMoVsZkg7BKG6
AaaUDQn7qBK9iB+z+ZisPVRFjegL/dp2DVoZBYyd0eK+dnJiAiEpEt/o7X/kw4iQY6o2fwuV1+Wv
GPAD436WQNfRAbmjEYY4FByli4pcXBQnkvgBZTP6M2z8cC+Oe09+wXWWSAK6GzJkVF0yAwssUFmP
l4SN4e4/tltToDsccpQsu5cH/qa58gXs9DSSySy6s1orAS3Gr2h31XjmRE/fK0fLz290Jt+6Jb+G
zm6qYr6gKze/EDKZVtZCj9vEDnw55A7dXl6gKxjk4T+hAk3laqwlyMNmdIFACrWm3Hq37/o1+fh3
npfsAAY02JWW/uEoaCPzccP9QozPwh8vod3j6ERLBlNnpRv3CWARICXtuXXKVyfEQbTbuEhq2Dbi
ir8f86bl7wN/X2BvdX4IYJT82iHG0kCKAirTtsrSILpYSq+wZJMLPSujpOzDI14UjC9h7WpbNI3T
Hw3nM1q1sxOx06bazzhm9f2dOMKxFsFFB26F0MmXPbBb1DC8ggAmZddEdXYU0qBmzaFe7VrMCNAe
RM/ZBmLZHmHJgPkqEC0eHPgbC2AD4TxfE+BS45FHUATGUUqkQg7NN1byxJYy5bi35J9og2oejRc1
2YuiWmwpr3e6x94KTgmfnwfWuidl2FfXMGqbdSgj/6Hor6PQaKVZ9SM0QgQh7KJiFyEv06330jK+
ZCmcwICp1f9um1voUTkdCk2dAiu3oorlwcrQpHBHQTdebD72aJT43PaRtzML9fpPqSz7zou/rqyP
qHjvwkfmx9+mHWiVeOV8jgsnoSyCJ1QQUO9fkd8zn5dXdrjZLhXlp2TtsWG1EnM8BL9X85eCp5az
BFpNDDE9rn/5SbxIl7zARDSYIuPZpNuJUj1ndqEMxayf5qsj+CF+GA3bbP6YqAVpZ7GCFoUksbjJ
AuVj65hQmkp3sDYcuvC7Vt9r2l5s2o+SBQPKnk+Lf4fA5FA0Fp7VnKIi+GP/S/C8Wd3T8LofPFyc
ycc7pmUn9fgmqTzQC32g7afiwI11SyiEFlyHR3By6VtLTbNNNkOHj/vebuQI8atbNSyOSlmftKjN
fuMl9FwCjEtW3oX7I2k2hjepYZ3skyahbQ76NY07S5qMwU809iMEF9WjRGpKj5KAlWDYFGu60Rjh
0OFJdtywJUdvkS26whcD4ry9nHZXV8QVaTtUoeUIqAizsSRpwtvkd32HUE7Dkg56FX4GZBIrg01e
6UaElELg2BsbT0l97s9A8R3mNQArV/IB9+JMUl5ehcnPD+C/A7BUxlvXy5Mh3p/X0ekdc2sDwOLL
jPcA/Wd1ZmJowZu0DcI4GRW/9xdILf+f/GJRKUYx5tgRjOvtSvDntsBnXrxCj4FTngNjtPx0QPo3
ZCa4M8qS8611QgxI4ssQxnyOGcztXAKifRkI7h3HKbx/QgORJj1dSiqQqbSvsY6/tqHzo9/pKBJZ
1hmC62XHwBzDOX5afn1WF4Fp3UGzxW1U6Qz0EhQsfuoGNmi1Eba7Moc+3deYFrbXipuUhPXNiIF2
heg5Y+sYmkgEyKL94APJbwHGpQvSV+k7L9wi0PBUXOfW5ErzfmrwPm0UHTrMbsW6Z4BeYV7T/36n
86Td5cXQVSbO1QlZCwpYeGL1mx9KymV2CXkZHRe0IBOaSauyE2kZHLG3d5M1SMwd9Oui1olPHE+W
8lLAN9zqShQwkP8YwvI1rP9mb80m7vhdU9MRg+PQVKd6avIsShdy/41Q2/uRMqkD7QFfZyjQPYK+
RHxqZ6aENmrHmmmokXaX73dMpmjxCh4g8fO8hOwdaffKzCsl2E1T1f+6jnmG0xdywR0o4dIt6oVG
88Xfr2a50u6bud7MwqMWDLXYFl3Ce84B2IZl6yMTDUYXkxJrD3RQwwEKPP27PHTurGKuTbLQxsiG
3l8KJlRpTn7zB2SXkp0K07L+r3fFWaMYudCpJ3AtEvqTCwe7QvgGWSZYMvCO9MgF+F0nofuO24Dj
s9iLc9i/Zmo7Z5PcSnU0lOdGVCxSSN45FhlcnaPI2Js9a0RhGiE2mMcI51E8w3cGew4Wd1vpaQDI
I6+cdgFL8R0nXcNCDe+T097wk8Xq7q/KyHOtSGPOMHYHECrNm0nEZR9edjb9BeqPKp2xMAFXR8gp
l+LkWuQgW7gofKZD7ImYwbAYRnyEGDidcBJJKD8ohwIK3vwarReqYh4h0Pb39G8GdGD2JWCiOz0/
suqthnjHfBKqciNQ9AV9onwivoFZ/naC0yP+iW2I6tRfHOV0CYs1J6KvtMDMO/DVG8NKSh66SeHC
Jehv0sfjIRp2eaOGNT8zXp/ex2IAZSJ0YM0+jxzEP67POggRMhdjByx7apMSL11lUvomVfjzWuxk
EB2oR4+LdRsQOR70WDFviNGsP5AxB4vt/EkHKt4zrC9plsrwRfaa5z0bWfLvJUFKD95oTlLjlL9G
mLa3GT/810P3vFa0Ag9XS9LCTi/x52P6pZgyAjFjQ1K27dYs0iurgdowl42gcVwHnW/dztroNujp
iR75VecpwTtw6qTUStBbxlrFDt9bDRYXJr9k/Ky0eVhbeMUfQ/4vf3bZZSCRtOTh/BQGKplqH+r1
i3ejYVARkNHN7QKBOW9vkQYKLnzC4L4JvtmjHhFhquLMP84fY8Fio/X5wU46/kbUxpUg82HnJM32
8NxUhqecFyuYF+mGe8JACc1vrSE1LJyaLjXqQp04JC8sxTcqGyKnMcCoUkIJPFQNdBHQoBzjuhTm
zfNUGoAL8l+OgMTXYZO3fINozJh/rVlGaxMblrtOuHlWzE5IKnleaW5TqmyeK0Qj5CVYwpTxMmbl
l3/J/OVxktKeAuYwCFr+5aZI0GQg5yUmD5XIkjfIF83eI4on5o38jmm7X2dqY+hbdisw3Uvdz9S9
0jfZ+8QR4e2IwUBV2qWGPo326JvfPPlxYqyRg/C54/tx/JX66Qy47dhb3qK5L8Ch+dQzU4fMdDAv
DAvu1IBLFsnv9LAHoM+ZOfH7PuraUFXO9lit9SB/N8NinOVPWcD/l6d48UrcofrIUGvbq1BtYvo9
+gx37WJg47+82NXJoShrZxm3Bt47GKLZThkMS33LrTMRSzQeMOn6i/hgHdMr4bE0JfoPHi+pxv68
a1P07oGpwwTp0C/yPFyOuPkrGJq+DqcDfe86T8PNLoToOp9TPb+STJDFxDuzBy6fNXyeREQzKJK/
NMO6KAH11fvCsVjFWteT1YcbgrEDWL3ZCSddwLZYFvyVtdrF2Y81ObqL/4rmK1P0L8OUQTAwApxW
k1/R3rWVvVvtDUpwERIJish+KJVd79I1/oyOZvNsBkmrpSgHa0zNrJvnNZwKGfeO8raiy9jHKYE7
6LbM/pHE5EFIHI5SLTgoY1QDgUmKFn7JtDmv6n9HIQXNdcC0sjiDdeebD64hCO0HWFhJmArtjjMi
yBNwhwtN93eFXU/4MU0wW6cK5h8AKXi5bQ2WU7K+LdS5tccTH5l+KlLunz4xDwdItFQG2hVb/Hmb
zHOUaafwk8ra0YrxvAWHhRBBH9cSQ7HZXtkMXzF8Ya9CZN38AY+/LP/En8nVEiEcuHlEzPynQBzH
1fkhvcD+QhBAz5EHVcR9LZqGL9cddxHMNsSH4i0wooEsrvhK+npFDoAsHD7lpYxCoI9lHTw45JzZ
EpiaUwo8cSgI1XU5yyySDUzwIR80nzD4z5CrzclLFmGDti6tCftdZg486PVwnBSNXKhdE7qznSpf
/amDKOd9wTjVtyD+w4I477LPL6Ienwuayk3GWOrI/xipYD399N8YTNmXPkn9fWw2WEvnjLoAfWvQ
smgvedI9mLNGxrU0ceqHbe/RelzhWEzWOOU9Jpu71qcIYPcnfS65uIpRJJtWnbMIiwuR9xFhuhhy
lXEtRivYUyNrTzi4ufjDOMjztNVsN1ONrsg5y+pv4IVFIeyzZHRLXJeKdz44F4eNIqw+reada4I+
1UkxQfBSgErdWy33fAjfsp9FKJ+Emdk0NN+LS1Fw2mZVMq2SmVgajK8VPNTSE2txWCLHeDW6mUBZ
jCaZ3HfcpRvQIT2cUVQPYO94B+bnEfNtvWQ2Fqu0FrWITobo28/4LsMvAcGqbS89fpVJ4a4VXCWP
weDdaEvGkQLqUPMA4tYDs9Dw6gfpQWm0mlnldoeT2MqmH/PrucdORvnJJTzNjtWNF9WkOU8F0PVm
xKS9s+2hDUW7p6kt4wJOiYaSJaqVdpYT11yIrkoNHTV/x5TTZNuN2mkBBdl1zrMQ37FSFLiOITcN
oS7ecCTnK/FAs1MqDo+nAAkokOfVa/Ezj3tGqNa6i6qEew/vXw3Dv9MJbaNb7Dl+a5F534VALRWz
+QXOaZ8roZO6JOykDOOWrQcEuVCJBzcC+iV/HUyP4gTb+SecoNnLWI0nFkrZ7d2c796hs0VE82Sr
sfLC8L5BiTjLw3msAp2b0twiPD1nuWs+PY3//I9DTJgLyZmzSCAmzhpzRud4K+kHkRGa91qhbvQj
xR+2UOELFJ9zV70iP2tmekNQcanPc43y88DUN8d5cp8IazSxPWLyJkEfY8H9aEjyMFmoKM1TMDaG
ezHkKzDoPjiYanmjIIjGl+Pb/tf7OH1X/avzTpEt2ciXdEKDTyidzNHE5XUg1f6qyJ3aopUpvpyI
tFBPeytylZa9V0hfWo1noCm0LFjdNx5mMmMe0GohRclcghiEG419wmR8kRaiWMutt6k1FUnDf0Gl
qXDhj1/WHHgpp49DhlTgm5otrbASLERfejnxdP0p1PR7NTAmGhBhKWRANiN9pnMfuRoPK3Q5YqtZ
p9AD64j1D9v2vWIDXJ/wDpJ5zOAEzHlio7G8YOZPB2d0pT+Ec3WzH9rhPevGqivw4BH++S3+8OBc
QbDbo7Pek1hEQr1a3M5V/XT37l/a7G/VixqXvr+cj/FQqJJcv5gJwvunElDCS08U9HSaM2Se4fNI
/Ba8E3R4VctForopxlpBxxnqFql3ZiBOYY/Kg3I/fH7nNZHXBD8+AyvpHsNU7NCxyQP8cqDYVT1u
IQxk1qG6SP2u37usmBgcbPehMnKX800iiJsiL1clYBPJPgmFp7UmOgnuOIXb1Xwhaxmx3FQOe6kt
NGxu+7z27WNkw4NoM3um+vUrIlpzS/V6MJZ5cEnc82wPCiQRhaV2Q6D5HiFaD3izdhO5lReZlue6
GPkkonoRHvqY4JEfdozvRrsnKued+ilI9BKrjw0WQ6fV+mmngnAFgUZ9JmdWodrRTimyBeGsb1Z+
XaCsope/7Mi/GGNZipSEFVpZRV5CzTQOfmbIDS3/ZM9TOkcp4UiY++6w3NoylHzPM8VWaeAZbThV
7+F0NnmYsnyMeiV2CAfT4YRI2+BCcpMwb03GKVkCpAMDEEuCO4i7j6RI4JyrRY0rBjLR0mBj1AfJ
x0uep824yjqfLP5yfygrC0pvGsVnKHr9T0MfyoACRqsVduA/aElZLMELCM8pwbXYV8EuPegvf9A/
HTT0R703gFAzq8Ycippk0MWqd61BWIPSsynTRIAEyXd8G1/7XSEdF98Gp/S4/YERWUs3izRjNWcj
1YEp/RmSmBSRloCNObZ4u762xWDeyErmnDNd0NqybXCZUDM6TE4qZ8mJG/z18SuS7CJRpwCuLE2G
jN6SmtERydaKoNmdVQWyfIiKX+1pF1j2tT3jeoAtexrNzpqOzq/swDQ0l2KBX/1D1bVD3V1RGrCs
gbBIYqidq66IlassDwGGF40Prf3arZsYqz4QlQVdxEznIIXZKh4adg1BuYLvDFoIiU/N/jC8KAzB
OqyJxDPGHahoSqAviZ2WvgPWxQKJuN4dJE7xoTprx4xx1/BNCfE5gmgdiy5tRCX23vfns4WEfT7+
c6HXiMTUfGby1esm3nAhQ7zWc0od8sx2CiR9gn8MauuEOMwZe/ZA8VzlSTlK64Py7RWEAeoaLFuY
QcIH6aj3oyzzKA4cavHxJFfWC1eVCwxSs/iaiz0SUBKEX72CQeQeI6nM6BP/HwvupsuvpGR4Upq5
9cAyE7Y0ebfDXiDQW0j6RQSj7PmvPKQu0oRBPjBLzMB99q2Dve3q8jUsT9Lq0MREZ7YMS9vgRdaA
Su8phxMT2z0jYW+oLLI7g9P4jphJH0oEMUd2ALV7e2aADVMuxVS5Gg9mI5xKeDP9CpFUYbBpEpLi
bYRX9VLg31a+kRqJNJFrWYSQTh3qasODeUvpfPFbMiYhzydqU+B/l42aVgbB+RWYRl6cgWfM0hXY
WIH5fe0sIIT8UxJ6sRfF3hxwaQeX7ay54G1OaMkIPLmJW9G7HG5zNqpEWI/WQkp2ItJKA6KOyka3
fzTGqskdL4j08TcuRcOXY9Vn9RWTlAcBXbJ7B2bABuPocAiupmOEPOmvZWppRHuDF1NJyypmpkf3
EV7YkWA3tGhqsBLg0O5s8hFCWOlG363r8zZGvsTTslj7gB6se/aQtV1fHeK2nO96S/Ckf2wJx9kR
8l49hvGZHIvlqG02KfbdmQ/EYkkspoIHjKcV5MC4/JWc/5oRywC9SM8G0/77OhzDAbE1zY6sDo5C
wsyZ0cQM714pL6mEZV9mMsYcydt3kNs5EvzlYu34wD5Yjn06RKnJ2Z6NdXA33QGfZhXCcGZs2FEj
p5CmjbbFtVzkdJVL9vHgjvzYYaRIoYDyMGw78fqJYrRjR1ST8T1WMBdXMPPKV/nym3zrDQ8JAW+t
7qAdqKnlQFJBdhSOKwDoBV0nZPueamy7f4z5hSI/l6tXQKPuta8Q4i17EoDg2BJmWO1aFYszHguj
FOqB/7FRrwaSHXwEFvDcPvOsLAqh8JfOeqv/PJqnNUeGgOwXygd6GBwNOpnJuuppIvgsRVDj4gNJ
z6do2J9L47RO4p7uDCAVE6VYSqKD2GvWiXHp3GWoQbiiZH/pWdSjORkoyifHfCY270dWZd00nxq4
3OEDguacAsD7n9/vaCJAf/X4efBf1Kz0PIyzCGUb6h2WdTSftKq16N4kj/99fRFtdg90zkdjV/5i
qxjkmL3SgCyXeQ8MfzdYMgnp+hKHZuxtDpgwDJ9UwyLZFAADJx5NDozRd+72legq3WcQ11Prd5xF
qY2qOJReG4c/c07WAV0Y0dlkZVlMSMGzrgMqZfSUoe4022PRqoZqu5Akbi+NYh3us7oX7gWFowzC
odst1KQhoon5oqdrcO9Vcc3LChBKUfXnG7ID7ROFnsMH3g6RHZf3oLBBCP5u/JW0Zt+8OUSWsqQx
gxXkq/3S2VdxKYeJ4DNtiBIhNGY7ZYxl1BDR0UiD/0lC4ymkXv4u18EgQlQkmFSLYFxkFgvQGKRq
EwNoL4eU/VZxzhhLoCWj82qnIkW2UjpiFWI16n/Z2IUl07TuAeA5q9X9AMkGoy0MawhlpnAnOjpH
lKckz2QGqiBksYuTMlT0zFFUeSyYcBgKZuGB6HV7Wmf2EC4Daj/clK1p0Opad7d7pkT4EOQSTPWD
2Tn6KkHJUi+KlBB1hs7Fk9du6wbivIjE5m/fNI/O2BxhslVsNM5MvbI3kX9KWqcNZBS+iCMqq9LO
T6dnnPCtYqgWHBwBjBcmNdkuuFyDd6YQTGSxcZdm2K7soPu6fXUew7WRe1NidpWQwWOlrczXZCRp
NRdEVlXPy8IYgQH3bR7gms4ARGmXmlFTtsEvbEFcu7sSbloUV2g/t+Zl907CDeiNSQdxz5JXf1tx
UdTSUsRmD4dlGhBJCm5K179S3HUy1+GjhgzpnW8ZPnErqIMzpF1V3e4gEs9CGjaAqSks1ToIgaEG
vJktptxAhQ5Hr9eIWcBwPfiiGfr4Znpo6l9q+RC7IInux9yHeSxVImB8mt/95iK5UU6mJTdlv0Kb
u9nDEmZInCS+paQopsMRpOYjfh4hB7g/Qs4MpoDWYijZn+FSa5tnfMNlG6vpIj2jQtzNqPPVqEEd
aJZrZnjf64QRQK4wldgFUMtZB8tUCOTlywn4hhc1KDT9a+y4BdvF84wNRH7STojgKkWe9rP/yS6H
hCgmRzYC3TObyEOK7V+gy93zZdIxDHvR/KBy0ot7cTPJQTc87lb0E56FmvUZZYZKlZ+OJ7AbHgLp
BDDXidconkRCFXWAtoH86OwcVkSujxX0QUaKIka4U/6n2rASv/AB2qaubKy3xx35+mpNVt3KAxbJ
OddJjzKq61SJiHNVmzKE0e2n2qWUfQ0H7Pen9acFq2DdbefPph0PbzP75eTXeSmdelVd5GS4hV0g
BD86dp8TVLob7asSufJr3NBblqHFw1bIxKC1pZxfEHYq3uvOVKpr6Dle2rlc4o91p1UCxFyHlrZh
tuwNucv25nVEJg+bS49l9oLGFXzvSIOJTukFQhL7tMkUYX+jy9F8Hide94JDqqENaG3dGKjsNL2X
ZyrHzp2Fe0VrLnS/2ZJezNjCtau48ypy68z9/rfb0b/W4HdStkPf80bGQkRYJOykalNwsMSqh+k/
8/v/reMN1x40sDh9fVHTgd6gW2/4c0x/A56aaPi1pYON9AHSvPYf5FAbUfq1bos8EaoO+Ix4hO20
82WOSPINJmbqCOFDcxThnO+xF2yjNqogNF4oVZgjn+7fiejWpuCQBBjM3uVPNpg3jb4HgH6OH97g
MT+qBLrDfKlmPbyNUoepD1+a7QiaNg5ebRkqXUkugSkYYdu4nS6n4RQs1E4LqttIpPrXva4iUngB
ZslrlC1+v906pUH5WTllEZ4c/IyM9Xa+tFNgLDVIUhb34tqUlIHnQNEheRh90ynKmUEX8bb3osEf
spbWqoUCV29UQMMYJZ+If3ytUY9nmxrz9iWtLfo5EZuq2PDHKRsNy51LA4yhT8Q299oTcq2RAmMo
8KTGS4zrhIBE6SkdtEdHVD5VSQPC1rxw9z5/KcuY7gmtj8v6xv3ezEPL9WlZuxt10wfKf6boIVPf
+PkyxpYsQ+fCij8bHU9+j8FFwWhVtdZWyvEZSdh8aC1oRvLQ+39Mu8SYoiGWtEjBDYg6zrYchW7d
C8VUTiMnjpOjBMwOMnvao6FJxxV5FB8eQjl9926hc8f/vxB85sQWipzqVEC5QO+yVEc50FzTMC41
yHA0km71PpLJGst4HDwXnakK9tSYNP00AAoltU50Q0mQHcrzKMotiDkw3KwYq0SIG9ISA8CbM+19
9dRJJ/DAc3F4sBJevutZhsfl9mppfe+DH0kM1kS3Wr3gPbic29GjiRPdy1EuQgc5Pphz+1XUsQ68
dI0D+HYHrB3k5tzlxWnUbYFVLegSTwYJxMduV7MJ4aH0OX5uS+v/6EAfrTofXKwmxZfUs8sLRh2G
Vzh+oWS3/5hqtghcVOfsWg9HPo5+GoE3oDiFG+vnggn21uhEmAU+jLJOSmSI0L7Xea7J8No17jJb
ng73kJxJ6bSxItSmKaPGl22V+BQ65mosLmL1UG0n6s23aLhc5uEexdqjhoEcsLYvhLn63XIzkxg3
ZZba9lsOMaw4fMbhymdsscyVrAK3qRGzB19igzPD6jDTeQM8rt5ivYt+jKAWIg1+cGcJxkmcTXwx
6J3zREtRV/QCy/o50YDc67yUyh7tj1QdEIlN/NAdmV4nRS889AtayIhe3JcV5F6SRIxNptRgKMbE
gOqf0UeB9wTjmhvWoeT7Dy6gkpMF1pyZsUWXYICIUpRqGJd677Bq36WwdKkdeiCj7nnR5t3/wYPw
ySTYQE+lp8lG9KF5NKTqqu+h5WH+OLhx89ffAdFlyPKdc0g8z9eQf4n4oaG4VNYuntduXDf78uSU
+JePAF+TlfGKxrleGuEVHFTJf5Lko9PFeUJzAlAbc1dFnOXDysHMjrfpDzTKxRqJATyfGD5dZhRK
cRkz2ikQeIZ4mUvpRb9wR5gITW6y/eIx7iKdQ4/tBqrsmNQqUt6uBSkHwI7PZ8yI6lly+VaedNCl
4bE1ZkiJtO9Uwh66uCgCxlZcc8QF0YYVRw/SS468XX0fOx9txbTfK7mP6Ut3lwKqIuFDNGXMaH2m
FWUrBS+q0XmkaNunUaASbEkKwbVM+B/+BZpIgj6fa8j5rtm4FNrMMm5UtSk5dolt4WFeDvB9yomA
P+U5ZuwzQi4QMGD11J3xGo/Q+aQZhaqx7nqj+wk8eYI1Xnp4Vvbt1bxxXMYqTcw47ta+oAmzim78
KXosh9aFXocnwxHk5usA5HYfLXos8xe9e5iEjmq5bNuZtGWQkrGce3QhRmX6lYXBowaPey45Y+NJ
ScqKT2ib6UBd7QgkbXqzECCaWMKEgux7uwQ651m6GPuxzBbPwGLIdJ+aJ7ktpgNwsx3+65RAt62Q
l1WJfk9Qu6EKbgflZkEkImlJ+CHBm6xT23KjICUUjF7/uPJgIaOOEBw8C28675jKP2UAIp9FuVt4
vgaUBvEDqoXoU3Qt5Oymr8Hzl7Wdc/wz+rY0hb01Ugz83r2zYtjose5xsZhGcnYVt4m3cTupTa9/
AYpZ1b0Ti+AgQ3h9nW51KB/SmEEgeEZkke3Q/lcWYTMt3JmipRECBaYdbw3xjK65z0Ny+cgxJSEK
8GKWODE2989p4ChoVXl67jVPhB6NS9kr2BwdJ2ZLpepvhopAJPuF8bK0MXZ2/8uMSmrCVk4aRHNN
u53/lkTmSY1rs42dIIF+FrCSzWvSynVF0ljyDvYgp6PYxXUBJn8H30QVAjNpVs9ZbE0pQBGsLVuJ
Lz+wUz4+XIAphW7OhZRTa0QDAzz9p1/493gzpnMh8N4Ci2J/oXJGfxXxHRZYK6AUD+kaSO0GGDUn
pU+PwJHkIVPtZohNIvpgA4aKNWFFWY51ybddTGN76CkH/aDvgUJShSPwmEqq/f/D9tqa5fesLMK0
gmmJmV9ViLADljpeJq9okV6WSmfkMHAY7rkpIg2dhzEtr9LiCXPqFY8MWxlZ8T/lDVBHmlrOAclj
iYTQLqhANZLUKqQNRFPVbRX/UzZwSEdBXEmrArfBIp9qZNa/NEi3bA696dc9gcm0uVoUPJOISyep
AtjoTqUcbnFWu6POOC6bP4/Md9jAZqdrdBspem6i9Oy5C/VO28dWunAQGwdOauybKIcAeyMYPJ6N
g4vdKSRDe6bZmpZGt0237+A+VbgHxWqhArvMtcbPW1GIgqIPWY43XjsGqo2TduXj7pX3R+Cxz7ns
myPD8xcTq3TgxALgXMWh27OJqU20p/w/9Qz4ERXsQSwN3598CJm47jr9ZxdZFo18T5tsa0G8zJtQ
JSrQCsBQ4Z9gyMR18PAUvYdBotNCDLGOOfYN7ZW/NC2MC0xAVM+Y8BD7xS0ufbLcCmqGazvzg3EK
tGxzEAoeweJdHQpTwKSlpV6kqSBaSRIsBqVqLWaKAamV2bSjXBGwZYDaHvm5pfeWhlKqASsgLJa+
sMMB+5w4MyqRAa93sgtZs17OpTI6ynMNf0e1hCoQ11uj0PtYdU1Bp2SuE8m7VTXHpWy3qP0jUD+G
UkGIygUNwd+rs1TmbkouKUMyBGOmBhmgEtYnUybrvFKrxR6Q4uWG0T+3S17K+4nx9Pop7gshM0Ck
L3Vxukph6fcE0PCqlxpwAZrvm1oIFygpR3c9jmekxWIX6/ihH0UDIFlpQhgSOqnRfmirPfoKkMrH
/uOLnCI50T5vTaWkw3ZedbdWZ39nOaoSJQvnWH9pyqYKMXiDQJrIjc/dJ9Ilka410C9hlmJiQOx2
fPLmp56CDElN2CcgKFMvuv8NC0mfDXNUv3CETokw6OebqzQtXL8fXzSVgMqaaJ+77hqGPH16d7Cx
DU33Crfx+KCOS08H/g2Mf9pJij4J1gWBGYgIUDXeyzqhshht+t6ZP/w2iRRzpzsIMhfJmf3PYoSH
319P0uAVhwzYW7dixUR3Jy5j3cDzlJoW41zcjzBiAh18PnDUUbGYJPFgk/KNKUfifPM5sbOXtaGv
WhF5rEzc3jQlaK90MxE1j5+EvNAH+5x6JSQerr7xSND0XW4NMiAey5tJpG/91RoabJQGESs2r+um
VHx4EyFNYIVRRbx4L67aCm65XctKqZr4ig7sgx21BvPsMy53n08pYCV18LD1pr5MLJBDcRGrjxq2
FC+71bBshFVn8/1LHYSBBVOgtcqrSfKhbgw8wGa0KZyAusOHmN2xmapFZfa/Bj6w0t50bYSokvMA
LqqVgm3OGC7Qt9tA1jncEcq2xXOHKWu05ZVkPoSSQby8W/ji1jogA5/1AkNiWCtS8rl0tpPh8gcT
8GCt7c6V2bB9j1ojT+fjP7aogN2UF1iRgi2K/UsuA8fM8dWNjoULK0GZ+hgOCtdfuDyPLo/Z65Lf
dXuhWJwIwjH5d3y/OSeBTStwbkjYqno1P1QXh/lFzMEkzTlo9QF2Bxt0aFkDG+vihGPT0E8xK+Yp
kXxPttjj5HZ1hpeJv+8v8lq0SToC16r69BK+4osy5gpjzGw7Kg3MQjMre4zI/cBSEFKFa14XQOWi
yn0hz3+mUSREyRX9SBB9Ggl6xcVDyB+66bKny3p8m3ilEel6hr676mzdb4oITaumX98MOmzoL46e
ukZfbczKSkMj2baGiNe6Gw4NtryMfKSee37kbHf8OQQXVZwbr55ga0PZIenSZNaMGSs/wJVgLH1T
+ucF5CELPBpDsBHFw/4ZPcPQiIKhFdI23SsQ6jGf5CY7zBP9QEHy25hlyhn5DWuyA8+ivqXFJvEf
SMm3HsrpqOh+90rotYESVgosNwblWpDyn1VNGkGxflxO4xjGPWz8t9L+uta0WlZxI9hWs0g/88uz
lO8Q0e7eJ2rwpJok/qfXchRmrAS2eBQ5p0YePJzMeUPzbqfiot5RcMZwjS3ErMJ46W3NyuPp8IXq
Elp+cqeao/dwwbb1LQodYaZvMZwIo+SInC28pHZDXRx2xyqStQr0Eh5xMvu42g1eFPqFen4cvpQ8
zNhhkiKQ0G5Ydtf0LQC6OMuukoWX5nAbgV23mriSlIXQnd/M3e8zTEmE0l+l9vexYJyTsRkdpWs8
ILLdeiCnRbGNGhmPtugIoIZ/vyuRsJUkBygBkdDmIFGPbcL4HcdxsBk6pnbtQeDjngu12f/C0jaF
6PYG5EiwCbUTS7bmf20j8/CBRuO39F5vfMTnEHTIiBDGTJwiFgN6ngvryhQl1rlBlrYzQPb0iH0K
LKkWuRamVjSVe62qZrmF7SltUWwJJNszvf/NHi80WD59or5JsY3vkLMVloz3ue7+RtQy7poGtuFE
vlm59kEsZMzd9by2Tg8GrK9venR6Gm2DKU4ty/b2RJQlha+Xy8dlF6DcnE8ueViYrp0E/1tJWjDY
I7u3X3xFKtUiLFSg0bJLHkebC/hHgby8Nc2n0p8QtVPVtC+N5J1JB1MVZqbz+nBGZvrL9GY/B6w2
t8MoquB5D8a+G+Un0Q0sj6Tp7yV2ihd6tdZJa8tj0KwnEBwuOocGTkuR5nWsyDGgTxa+It09s0K9
hdlKBTvG6SAOqI4UDC70yT5HQ4V2OmRCCBeurfkiH2J/vk9vRJCJS4V3WjjK0f/GTX4xNRDddjC1
WVspjlyefrktTlfeCtZWMJAjuZkncYSteE4g8WGH7wd3o2LpUnFMQHiHA2FZ1doIi31ZrZdc8/8E
+ygZgNhz8bPhsxKCTO/514t1PFbd4SwR1cgV0D2g8aMB/Qoei8xnrdzgupB+gruxh8EHsVyEpml6
Hmy5yy85dqQv92tZDyIQo5+5BT2D4gj1iXaLuLu0k7NALZTi7LMbc3zr83yL1Xua2n3M1O94aXUA
Q4Og9ImJ37t39c2fUcV+q9aevvhWa/NDabqFp0Zo6El1zfhdEjB4vUzRXEEFoNLP1duPj3O8YuwY
emS9M+gI/7SIRR2wTFZXsOrSwwoTYaRRV1r0VSo71eFT1biH6i2PjmlMmT7MbObiQxjYnzefFVRn
OrqEW5PvYura6xhrXnVF7Tc4BeXFZdO3g3wjGA4ZJ1Is/lxpZWCoSNLWToW5hyRLNAVq3bCMp6mM
KGFIU0ougB10T4Y7NJhnwe45HWefc9pZwBRfwvWxUqaKCuzVtA+6r+PUJPBRLWtLTaFV9t0eyMPg
R+y6wOSv/SLmUmi52VOn+DKGlIjEkzlbgx6ayOw4N08WtUZLkxXMwqwzCwN+/JlI9IzR5bw70Qr5
dT/WmfD42E6FW8E6IjRcjZuvMBXfTy841w/VwOhbebu5p4Gvz4BZtweo1E0xUs63Cd2TFiuadKjq
/3zGtT965rLuvklUwxfjqeofTEVpr4GfPhifUlgz66sOND6e2mC4wpUh+r/VFd19mzjO9hDMULbu
klpcMb/nC2xSe41Wl4fNefN+ZoZMUszdjmytNWlivj1+XLRIBzE2wQoY7bMGdq6IZOOp5LG4givR
lWFeORGWqw3RTNH5TAuOzC46twn2hVKzJXLGltCj6hTEf51pq1htDKIsM0fHyHDQqnU2g+YnK+jT
Cl3HLNwJFdrLjs6IQpE805z5JB0HRhTxS6qQ4ckaaKHGTv/sRN0S5ooBtUAeiWjlm1x/Rn6wEXvt
WNQJ5ZhMrOvVEJX+v4W39k5L8O8/GK1PiMDasexzpAI8zApYUP4mZC37HJ1/NUUQKRYC3OMVaaSQ
Eusx+DqKBd/fNhM4AiLd6VVl0k9tyIcVBit3l2BLSQ8aDt1DRgA0b+pEjl04SZ81Q1I5/x+K2OeV
0CahsIL249zb9X1l4J4A/vKgM4nN5N9B55RW89j9HNvPnKz6ypWtjf650y2UuD6ltMq6AIf6DM+H
/4H2AYOwvKnl5pm72tyGBGgdXwm7Jgb2z+xlt9BaqN1cwA8Y+KLKW27k1nTFYI4dnbBVLj3Eroog
1mKlr7Q9UlGPz7PTrx29Z+hPXbEPdMV6X8jp+NHCwSOZI/NTUgLgy/3AZPe0NWo3gssPInK4esTa
MjS/ZYiAOuSQizLY26wQMV5irR4fAJmmQLSUA3eSIlYloVUMJtL289ZzZjnCNoygbG0p38gK6V0K
nbIen0gERB8qRznc/cEKUYPDSzqsJGK0hVnlhMnySi+2JgW8S2TnWzwk1lIjQhpBMCiI5pEBOa56
uqp8acur2VBa++3wfRlVp2OH586E1b2d7QkUc9ehZgBX1cho3Jy1sOKT6zVeFhlzof8/cG1LTWAm
nYePqAukZpFwAkAeVbxS3k2BvcFKnh0/o/8a/7CGLMOelqbcYoF+jNz0FIpIB7EnIrWta0GUXgzT
YDkMcITEc64SqRmCjzEnuxa5oszCIAC66W0/G4VQpHwtRFFiUCWQd7wpG8UITT8LA1nPXcKiiOBF
zaLyGfM9TY9x3ZaXTHMPu9VTARKsCYYlWZV5JpBoM7SKUw03WDmPoM1PiAwsg8xv4BuUaFZlpCSr
R0oDH7mCbVYpXsn9nu5xWX747/sGddj6iOT6pT4SJNcNwkpA2NpaDXjs91WK/dAV3E5vGiAL71mW
FgE/ClhBoGG8820wdBJhK2IAKU1QJelecJCr6roDJhcxfZw8H93pHxftYOGb6tJmxGU70NPWoNLZ
87KiGf7zscfg944D6FEdEN01h0eA59lfZPUEa/F1c3v17n2JTt/lzu2UfvBfNvtD77S2Og6OyKCQ
OUG1wjX1tptCqvIe8xKiPzlDpbPGR2V6kjca5yImWSiHY1SkZ9cW/aOYN+EaIMreUwrFdonPFgcw
RBNoKatJGarUB+G5BbwVPYDDUx7YiT3sDCC35xXU/7Obi6/bJRI4ZyRUGKSJcAF4AMINJNgSn4Sv
kyIbdQuCgYa2I8opvhN9guaRYCt4Viuco/Ltjx9VnKz1/W2pYwkqPXL0BRryrJSffjOjBvi+rZ2w
SNOr4GJiRG5/Otwl9GdinM/Hv3rqOF/qYP+h1W+5R4TZfBXJuEN9OG1z7vMuSPDw1maApUn1+775
HfKXPOpMNDhbjKfcsiBxDPxD0FfPgGy5k/DRR8jIdcVYQEOm7YhBTTbeJgnb6CseTG30kURFXXrE
gdmG/siu/NGSCWOtOCHxq73zF3FbnWOqqPmLVJsFKFHH2+Ps8AdARpV+0IhAB10lDSUFhAkXYwWs
uebhGGVxonOXLmrZX1IFYdLVJ5i4KbCokvll98yYDRVI3gopKCmmcwoamoXRc9Faz2GNk0ShzgW0
Ra0MSyFg61La9UoG/zkn2aZzZoFIDIcUDjcgxKitDvkTe/h6jvJXZ91medBvHf0wGRPJYT55oXVQ
lJfdd9j7w6O1hYIVhcGZCz5N4ozesws4QyX4mT/Mqn3chDu7tTT4QxIc/GjT6rFWAFU8z+BRWfHa
90o1Z7qsT269W64oznGDZJxv6vwwp784ZLp21wkHJwUyBYiQaPAk/Ut3ejtR/AhR6QEIhVyGaECG
+CEI/WnVHYFOygm/NAFluj6jqQ7edszSUb1A1oi90AyChD8/Xp2LVmMzLPItP1mheOgrmW62oUE5
9Zi7oujqyqzTtxU+4ZVVZt9qqcKTYXI6574pE8ciF9/cZv5kJsxBWO1Q3hk+cH2jr/SDKXnh4apq
MdaFFqIOpOIX/YKfDjpK//iEAs9qkfEATN7MO7VKQ646ncW84SQscGRVQviZD7yXX4NVUCx1qvll
sR3FI0jCUK7YYFlIADfW/ph7zyRV/4YLs0q+JyAhFF+bpY6jAHwsKcMktJEO22Qt7vRjTaqt3Lr7
BGrgtWk2nz4H5H3/iXJvh8wah/yJe1OsmZhx5iN1zhT6H7CJ6SZglqJQQ2WLjcbpoAjxeavkqgYC
Wzx67bprmQSEc5wKlEbC3LulP+NSAnzvdnc4EqmbKCAAqHJ1Nxn9KMuJoItdVisBxOqsr2fpBeqD
P5J5CEgVRZvzUtK7oC1t+zNPDbLGFP/Dz9/t7igJ8afhri2TxTxCwSTnmkbY4J1oA6J3W6NXB3cn
LTgT4xy5i/paGJZ7M8Udrmqtu4mc5vtbcVB/vOQpwSYKXg9htHoFnLTWVxBwBmZPthIUMHu40gDH
O9pevBcfF3cpSLW2c95pUrvqwr4OrTlmiUXLr3yu/J/b1xRhtykKvP6Xra/NeQ1t2+ayNgAC40c6
NuZUwUNno/KClO337CVyuUyLVD1UmtpWEP8WvJGp4bwo3kvsXPvxTI9Yc/cQpUdPqQ50F87mvnvh
JPcvguI0vw7v3AiMVdA2uSP7/7fHcemLTJH7grob5WKFY0DJRDOO735H+6Pb07qnkPoi8Cd0GG9/
DM8bk9YZ1YjDK9Okh4ZQxhkRNz9U9koTuEcQ63+/RElhNRuOpFv2T60mb08JdM67yGsqapMijSLI
LO+9w58WrV75pGwaZaWdyFPqXa7/OZgVuuV7YbvRIg4Lz0D3cdzYGFBWwhB/sLmmFVSnjh+Ze730
KtnStMKSiCcPLPaAFcIdxFEVI5NVAXL6aZ+UtthA+bYwgIDZXkZRqyVM3YpqagzNsnV51oSXbQSU
uKV5gCPVG6gWo/AIR8XDKv+eP6KLdaN/BiD6wAx9AKsaNDmN5waFV8s0MrrV+r9MHifq3oU1l83M
z7pf0m+j1AFzjTsUcCoKzINdNxb6b+LOSQs/1jF7nHTZ+CdJmFIIPYurqyRYSFj3Fu22KSgSWZs/
bbpXO21/wWps0a4jHGtJm3LhAv/6ib/dPBHY4pGgzlNI6Pl5GpAhK8p8d2HewdLbr7kTINTZlO/7
fvfEJZ4EhS5t8x1osUQcAdT3hZ6z5L6G1k5vP2GkhZ+0t73bJsEfskb0C+WonLUfxjvDRJrQu/xg
cBNM/daxILC2smnkLSStgozVeX/ClPPgqTmcTHUJZzZgW+wrPlufIX8PN6nWfLrG0klk17LMOGOO
DpVbjEIDb62OYAiHiFDXgkJE7eEdNFlbcms20OndzvkvA4UiQnhwVdzIFsIIz+ioNRkhvFKpY6KK
0SU94frWkz+y40mVC2Xj+2zUXJTvPXt9j2+upcqhc6ja9q4XEoWXaFWF+0BTHluKV0Pq77ieE5uA
IFFNftOBaoFdTUdyA0ZRx5Pqqq/SRUrjcfRerwq/RqOj9Ky9U95sPVJ9IgIT4F4TqtzXFmSXOwn6
y+JP330N6G0cLTrfq2mftR0LMnLP+OACED3uKT2SZgRnl30QTdirMr7+Yt/hsgqLrippt+uxLko9
fro9v9eMHebSmchpZ9Fy/GrQE9XK2q3S3nd+NFMsZE0O2DekUAzrpix9qNZQXEQwR2DGKcFbDlOQ
oN+8qcyMdikg8fhCmL31dUVjA0vXNCUY6k82NS0huQcxo/n9Mwz3SuMO88FwkKwnqNVB3h1SAe4S
Gyyf28WforjgFp6rTRveap0iILkeDk5S4rX/XAWCpIHYCSng4czYPuzFNi6c3uI4oNW9tnuEyXtQ
mVwu/zRNvTfBw0IBl4VQXw0BG1QrtVCutjjDSua63DO7CIRZTuqfNTmkvw8W9+D6JaekQZbLpHYF
tzGmeY2Ya9PVMsDH8Wyxv2+3a0pOh/pMIU5MWDB0mek5mfSEGd+v6xNF2QwhUry5ipRbdixynK5S
IElb9/Ya6oDVt28by1BznLxNtLjcW/L8mlO/8LmGOL5MKgBFdprSo4jWj4V3ga7eiHlErLWzLhyd
genwHrG16ql94IlP/1exLm2x9a0l0w7VGLl3/0FAYgUNBcA9DViyfkiVMfgbaljpfu3tAWqSiktf
clqWExihx8+zIlP+pAc6IlvdYRazh0MBisQbOqFCJ3gBPWJXsoHMCLEKzqp9FwvUiPMO4c7MlapD
MuwmghWdaVQ07USf8og6VSv0wJlLXXcKFOqbYYJk/ejYU8P60pEMFWXVBxHhdQUXEuhdUorIjEYN
koWAExdYADJQok8GKGvcL64LrFOf8C4tMVclMKPboYwFRN61V0ngczJkKgJWk0O5UycRrM3Iue6i
Omnrfc0adCnSODGqKE1e28fiBhIA/j79P02S2hV6/dD5nIKrtx/znx2pUtJc6572Ex7rzji68eVj
skhQMkJpVqwrGnTwBxvIad3wCILCKVio+9Fojr3f72dd2NhfuSoWa5ewdjIFMG9wHr8hQgPtZigM
dN0yjAWBem4e3/C1JEEP/XRuJTzuzgOggl6Km2Mnm+ZmQs99XvWhDdEaXapg8rNw6ARxqo+tCdTc
paeFVa7R9yEzW+XvtnjeZxc+1BgiV+iUSTKTb4RsHae/91uknIJX4wrcBOXwBEWoNSMxSvDcR3CI
m5/wbKDEP/GaVvrQGNw3GwV+bDjHeYEyczcastjD8Rqf7Xieo2Pk3/XE1gAwFTjh2YDJ+k04U5yv
H9h6BLMC5l9ly30V78KJGzpVK5nlT4MlDICfJ4p179cDc44YWGX1BZlfbcLrSQfHKszkM+JFqt1e
jwRdZTZuBelShwwULpYstDL03PNVCn2hNGbA8briYKyovN1DGCjVchxT7UdknWR9pi5QmEDPo0vf
mzWSHVhBbfb/ovAW785i3RucwBgXe1vWdrvYtsI2hv5FLjoMoVu6BHFMXyRlYg3PwVfNdCHrn+Pm
sdQosefzAOmUoE+NUgmGsvFWSvhtd9pI4YjnSYBaZsYKVJPlGA7zL9deMMm3YyrMxXXjLSzr0b2a
9rl9tY4JSrgAg4ONpvQYCQUf3H3UdkNQcz7sXQqMn/iLb98EOPK1aar+flcDQTMVIHmuS91bQCwV
S15SBdLqpRQG4pOIGcP/CRYNUSwrNqd+9WpySVJA9JGkl2dEXT8Mn/H4MrBou2JdSszOvGPVgGfE
G8m/M6OPuC0Ft5hcN2S0oTE3GIrP8uOiUPAsVBjhHJbumGnk+OxUUELNsku2NfK6yCqs34MBAlId
jin9Fm6X2mIlmwd9Bsf/RhNb8AhHFg24U6UthKYIX5HmxafO8bU5RRl+aYVfl2bxPJH9QL+oWofO
c1z0du0ZwxiHKo12dGNP60qvby+qARfwFqKzgqa5wdni9a8QkRErKrhhTW6TbhG7N009XPldEDay
itDER4wT7NNdReHb9Bb2iootBodUzTnvUi73+KTunNR+NlHwsFlfwAIfxzGBnbyi3QGh5gi0+vNm
cg1s2dKBrZ8f0g7bCp2a3ISX4TJHEaQPOX1fH1seoMifzjl2Wj5IJf1qo/V+0K0N6Px7TbtVS7zd
2DIlLObDMcs9xIV4uWthrhQlNb4Fb9KXyKothJaOOtxeXUIMNNb2OcAPs1W9i0UPhjItK9HJ5hD0
bmIBMSrQQYbFOUdaLYNmzMeEgcEWhlSeODDU0j+zydG8xLL1NOuKOiQxqwJeFCSyHU9nLEG2N2wc
pvA2NRx26lWEMuUnIzwObx4vdz88Eqwdi7F8Z20/tQEyiaPtSbSIB4n0LBJ8ZGYBJHIo7YwfuiTl
FrUdGaRyKBLNbP2oXeqvIPmQ/cFD3Qrv7CjcGIs1EtGlMrFOUbNpFdQq17bzVhLIsDx0m9Ptie2q
s5odeMBvwRZMNgIn/N3eL2QeYbtwD8vndKQRYETlYYkApJbW6JM/XE8IXPgz+OppSWlSK2XRVxgs
a+oEqEj35PmMm532dctWWFemOb6wY1W0qvcAxfqxLUEZWBtM1OxNNXi1utznzhDRsOcbZT2gNp54
PS4aEUMboVomvbxS6ao3K3L01b1dKSFuB0og4xaufnEehn0KDnA9PuFLcyOvVyCoSnVLv5DE5WUv
KrIL8kZJAFXQZZT8E9TdPY1kjcZfJaSHyIFgj/SNxmRy/mVSBvxUV2DfrQD0xUMHDuqqnVqZ/RM3
vFqgm1mNTpnyjiyZV4wz1UF1F89fdbeudiyosaTv7FeN+aCckOzH8YvyAFRMhZTgK+6PLIufNr/j
QCq1xBiyps0kMIypeR3Cg10vdQfu2NpDKYucaSN9IpGV7pmd6tPC3k6dTsCrPAo1LBdqL08OvsBp
rsbAi6J9/cXN+LqVrAXqlclA72ipkH4njiyPmIpj0ZOHl7cwdFY3T0jIcYyvD3pZ6AjL2RoCJpgC
2MrGNbC8btMuKrNgpNCo11Gicz0HrskOvPuWa3D0i7sEkvoo1UUquJvR/3KMzCVOQ3QGMAo14xRP
FRi123Tiu5XqyZOpdm4R5GEgJ1OkpeixtEjPkVoqXxUEqfyFThhnzrnMhOEmiEbbTpPzb+dskVQY
s7R0llWH8RGnVFzxn+Zx1iHtycfIxCbd3DsdTEUwG1rQYZQXULM3hBqH2Z119ScRsSqz4VWhJkiL
tfkHikLl4n0Ao4dUhUx8PuktENWXpi+Dsj7LwjLFActgRUNslATs7t04DPsPkAyhPT9ijAqqf/Ty
dP7zXlExcl8DDS7ohLRvfwxMTJ5nfrN0o5XqdRKWwsNBOAVDHw3YQGVkSMJYKiRTlvo5nfrI+Kbd
oenmlsueqQyKbMTbNSXWBE7DdIgg/3PAvHbqzqNwee2hy6KPVVE3fnYjvZkIGd2keOGGZbc+72V+
MCoPcdbHhcMCyN0tHwtk4S5R8+h4rzjP+FT2q3CXCRx8Ye4iFlW9hqKtaqaIqyu8PDam0bZtqtkS
Wa6/SUKtvwprY7jDKJrOOM3PT5qHfrMeMvp9aMMSGUPOWQqOUHOtBww2DscAC5K6eCcyW+kJRV7S
YJNHMdxN3SzZgPUiN4Y0FzLas4gGulSH7Rt1jWZnENCSTXnIDd1RTbgQXMO9KHZ6qe82NlC3GsOv
JaLvIlTs8XTHPcgo3WuLegQaKmBK/ZfEjZJ6Yv2hPtrQpFwcrpEvPi5SLJcKqnPOcDvK8lq1jK9X
k78TR2vHc2UbxcM6IWfg9/F+hU5xoAVI9ZEn+cuGcsdym9WlKLuLz8EBZQrlk/Hb4qY3i3mxqhfR
QMqV11J1pdt7GRfA1RM6Kv7P2oPMW/HZ+GkYQhSvrRaOp4wLaVFMR1+ulupBCdJTMIjoahVt1jlw
ycckjRn0OoNNTSwzz/AUtiW5ayxr/4CLDDXvG2mfiwwEFssVWLeGlL5T4Pvbw7fUjxyBl545U6i+
x0R8i+4UMkKsHhH5kL9u3bgDStx4AksXN+EXcPdRLTt0Ska81vYFK+peM/TkDp3DyuAq6o1pu911
f/AvhMCYXESKC/OpLuQpbxOShfbvtp0rs2/w3p1GvXikwCkPBO2fo3t1Siali5hMQqers1wjB90E
RAXbRvBCjJjMhtp5ZutBFyEQLawMePJUSktN1dobVWSwSB8GIdg9fhBXsJTKNkQBe5m8fHwkJDtf
U02n1BCN37XnTrKM1MU2yp/HTrWguj+GsmoYYUk6Wo19Sybl70da6PfglMiu5foeTw9eZSu4+zPn
U+XttIR8jIz4ASkniRAJ6DWJajJPRFn83Kew7+fOunGeG0R+LUeRWedhTavNgWHEjwR70eICNrbI
sfxuAqnrzHRwPxiBABur54Te1bPW0OCJE53QuCjTRrkY1lJKNZnUi3XSZ699rdXeEm4fdk/W0+x7
ylLpR6VNHNjeFrIlVJzg+VfNlmeZ9mJFrp1Cmsob4ANZSaNnmwkissBh2VEzUcQN8o3R3mkQwFGy
j6JlK1s2Bipb3PR9CbfgT0HgtZNHlpTXglUg/wRCGnrT3vrp7IxctLIpRThIRkqelKaryZYvaprB
EPDQTHJ+IWk7J3XgtT4O0NWLvvo+0TZ23X2pXW8UE6LhJ5FOVdjqTVPOyduIZgWT9wFymfKIRq4V
XJgvU2R/f9dTtRmRmwtmjJV53Y3n3+Q7YUU7lbI5m91+xdJMQpcALsOZIUQhotJVJc5LZhn0LEDL
ftvX0iJE3bXSLgL74OHbVzA8eDKy0ez6bYvpgj3MAUzsmQ5rVsoCYO5CQar9YpamfdCQdbLRb3FY
W66Vzpj+TKia2kokVv/3AYk0uuogch97pq81kKnxB/WPNKeNjZ9bmUVtc4/pmcuFQhMWorowAm3O
zwBWzEPSMrwA9DQQGOlKM0J5rmH93bjXA4sGTST1OsLGHWLiuJnHYcnA3LHifcCJODECJhQrfFAX
PO77sig5rEO1N9XVWyY7nLktGLph6g4CbqzJky7r2ZP80p3h6hs83ndUzTBU/U8+1YtEefpaI4uX
bGJqtUZYS01seAf5p8lPvKDQ0lfPFR6dkesjGA/9fPkwQISnbdCurljO0ZT/I3YlIm1MUJST3D8G
UrWw88qexy47PpU0JS9vhmt/fIEIxqcIzDJ34qd3KxYvoWN1k7IbMbd5D2OeK9PBmb0UX8z0XNUd
ITfDU+pWSnSm00ItGBk8Tek4q6V+qUSkiiYCOivNss7R5+qenHUSQ078A1qphJu+jFGd5GKe2kCH
/XqBEamNsvnJuJOttHZ5a5V96F1LL77MwWexTMYQeCA27HaNTLffOAprbU7Vn8j6bz9QRMtqzb4C
N68nRh3iUGFnLc6vOXhs6ss6oF9I50XnMBMQmcbBxI515kdtaLNJEjmInnyKxdy6vHCwrscZUDJi
IUGwxs5AAWu3eE8W7QXpaC8Jlsd/ahSDbH4V4JZRuRc/e2Yg3Wnd3Yeh+s+5sd4MZyTXoD3JRf8+
kf7gbi6bTwWrzWLFej+JcceFz72+EQ8WcdjP44XupSOFfFz9lse6TcrAzvI+Np/rRvzjszokJUkG
/qY+5Z1p8blV6FnvOxhBpeWer0O2K8Kasu4kLuI87jmcnB8zvYkpHJsl5TvPzayn36k7qS5JYL8P
SZsmX8BP9L8RjghhtEH900OpGP4l8Nl7tzOCqMaKIWf6Ki1+pWp1S9VuzW9EubloZE0uqJ4jl5Pv
0vVUKk3DlUp1bxy/z38ANVe7BlOoc8fIa1+t+znxvoQZhWbWWHQBgHlAb1Obbg+RO7P482aZIOLH
Lb7X8SKeRdN6ULiLgmHeo9MnNLR6HyZ863nk5+KyUWSwPJsF7wF7O20N/oe+K12RkY18LAufrrR/
jmA7PH1JilCZ57BPzZKEHq3BxV/jAFLCgdjFlAjWx1PEr1+mqvFujoApxlcuHvKcM7eXrnxRF4D5
76up2lq/uq9SZ1ZZs/q1t32+87w8BAwcccuXSI6BGupjMuL1pMLuHYHWi33Rt1UTez0PE4dlNOlV
LzswZ+HdhVbK9KHKjZ0AGyGbRF10qANsOPilcj8SzQzxKRSO16QtWT/hq+uR3/Y7liLHN7NqCAQi
zGzB9878zHHbzp3UzxEX4GYM7u+bu+g6WM6rmvJWE1qy8CpLX0Cq3KVm6drZPxi2kEOaf0y8+RYJ
tJlwutYW5J7TScBeh0cYQ1Kpqsry+hD1gNb1vWYTgCeDaBTjWNicrxfwa1XPX0aqROau/lRMPQhA
D7lJrJ1d+sB4aLgXgd8oWwnfwgrH3w0C2Z5um2bvPz/dMG18eJ359JXvVcZSX1d4lE0yZ71Uk3gk
4kRwoLgu+r+Cu6gpvd+HPSrkfrmfpVp8ZdUUH9Jf7jUl9e/L0CzzdhyVNRGSxZCH0f++xn7jRx+q
nJ3AWBPmH8B0hchQsjtZ2SFnzsURuTHT9NabFc+L4z5Esi4Hq9971AbOMr4irO/ZEPK+F/Azk7d2
B2Nv72eaAsX1waxPyHsR/+4/GhRs1tk/0jC+WgAB0jVeZoZqh1+yuZqcTsSph10Lu42nw5mYKpX0
KXXbZNPEP1i9Wf6BPsctioi5kycaVFfI3wl7B6gTnGcXkbIc5o4qZYh6+W1lfAR9s3YSpaVl1SYu
W4PWPkPxxRMnPFHxqwl3Csyf8lUXGYJfLdRDXGFOgT/RJanHvoMCLpdKiKBw/+ej3sp8klcj/ud7
HgATG5UCLq7brz9NpYwNpw5CDbXYsJjMG0jkSFMHRCuxYufkshoTitjGon+u8v2QYtCVv2DEwvJG
ft1ICg1gk2dwaogQZPLsaCwp+0ky8VAJzwkecKcOaqzq4BEuJQP1Msb4hxawqsA3qvtaCe4dgbRx
4BM++R0Du37F0pMTBk/HLq6pkDxwDIv6YCvnD8K2y+2SUedO3dBoMCpG4Z1d1KfpV595yEfO+dtn
arfcFY9mA87pQJqMhmJwG9bm/rAOq+ZBkH1ttrrnN/OlAA41a0YqVj2hlaIRJHzItcMqQWu2gKef
4V9xqzBLRdaPJWI4qfw0OgHVJbSOVCRgCcT4JzvCew63LceQJB2Udr19JJ0xjhwLN3ZbFsXFDWVy
8D0L5cGvFa/q4SMYUz56BKlCk1L9kucc6tQhLrpXon6x1aJrTJ8nnET6/uNOCCe39YgCfgu8owXW
QJVDTpw4TTHOZCUR1IzClKHAYzXqCI0Ix3MzSJHgnJDQyzSE937cbpNhLOx4cJ5ezGo1sr3eASOt
k7fftoQFJAKRYreuUP7yl8U95AND2h9un59fsUBoT12RF7s4u8DINE1886OHNrl3d8G2xFOhfN58
b4GALkBdIejPSlqb8e6VZYXTi4NpNKIAp6T47cJU0PQElGNgrb7S1CFSmGkADZ48WP44S+8oNUo1
e9x49ivFnvAjkmi9qqFLeL5iQKj2HiJzvSZ0chzEhDDXPgTN1hJWv4qAa4i9665vTT2P3lQZ/Nut
0z1+If8cyCtUBL2Furn2sFrNokQRINd3EAkSVpwx5Dt1lTPk2HTo5gxmzD0WZuK7ALfz3WXIPrwh
LlpNP9O51CsZWzEvFalGHBtwemgF+Tp9Qzl1ru8UzlAibzAiOSzoauhVapeR0It92jzZYxgLVLEw
TV5BS8JqBL1yeflAuqfvZq5/l+DL5RxPXg3Nv3d5nUyKFy466wY1BoeFJHels1KosajSFxD98dUD
XdgR1TKLzps6NkpxhQafq57pob1QfLsvnGaG3yMyKTTWdu6BVQ86/NW4W+Hm5AUEeLrNSGHI0qUs
yjpQED3G9TqF/8RDAVwwpPiuKF4JiFTceEshoRvvSVrF2tIpiMoJHRsf7RD03nRJocU4rtnT5uUm
8mDTwLdsI+iwx9w/C6hOigjZcZ3LXBt4EZ86p5WszObul/oQBPkalZZ6shaRU6qybYWzL52Y5klK
7labWA41/tlVTggT30eIrtxcPXkmotEAIjxCeqlW2b+UYGOSWey8QzAMrEjR+WGpUSiV7WumjH9U
w18aO0zL09qOvYPbUwHdMGdQs7DG5Dwd6fD3jTT/y+pllr3WPj7cKIjjc4UVmR95q1YDSVe1563w
dicSp4XbDzD3+4NkP7So+meD8ZkcCaeXyuw+50Sjq64x8DV2K3dBrHPjJXZiBnR8v5v6Z51eGUqw
nP4RBBZGfEz1CVDoLKHBAWGs3Zyl568bQIMnBkiHEm6Qo4nfCm5Mw+hzigpVmnj3Kz/oB11/tjC7
sSsKsjUA4y9yhVcL+lxhG1LkwT3KXpQp69j0oiMwg4K+Y86R++ZAEDLrCHItgt5VafpCLA95JzxV
3L+JDw2duu7lk7GHePFSDISQoiiK9zYt8w1Se6ARlSSSJUXTu46/mTb4D4VWaiEQFPc7eO8J8DyM
8oUZrqGUQsXG1M1Xd4AtmdLieknALWQ3GbK8jwpZKNn/Q/QLNkQU7BqDmuittt+380IfLEzlMX8U
kUWAP7OHJtmlOTZRn4qua/q8Sru9+CpsLVtJV37iURnBhdkKRMAPseJt/ckoEhSN0IOkiocWDTNb
su/XCb5uk8STp4uNUmqTwFRhLVe9K4bjbNtapCpBkap+6PLkIc0D1WoRWuukRYb4MFOPYAvnHw21
A1eM5yqY+sjfEv+hjgdW5YCPbgtky1eCEnwXKtPop60JVus/epFgfFhOG8nhRjpCI4JTG+NDvNBL
AeiRHnlJnRum+2PYyYQVGpYgn+yk3cR6aZ3WcL9S+qEoP9P12oRvLgZ4mFdH+DLR40Kj/eQ2LSSO
ceaj1u0JdPGQkrrCio3F6l+K6sCWY443LBdboGV3mP69VkZx48yzSMzyYPG4s52MgGdIXZ9u5DyE
eWBSf/X3MPJqXkwjQWx7244avYkhu4eIo8MFcnwNLL+NUNG8ElnuuMNDj37s/A08KyzY/+CWQe2b
Xb1nJcgqgwsN9aTItd1e/z0LjcgNXLOiNNGnk2bFnUfBX08kAgaj0HkuzUcuAI9uuhctBP2wOLzR
YeHfIx3e4CbPLpfMLbyVFpjA5DTn1DexcrqUQLKywv6FpppmCVgNkETKnfbjrABtccCQbLWiDI/s
mEMVnc0lXgwe+QmlsHD/gqJzImHPV3ITAEMsBmuuWKIIbEnhLuqyCVHtBHTgfWepokJENeIk1vH2
K6KLNMK3UJMsvjXWlNqon9vtUGI7Uq2iry8sQCpqUceRA4UY7RH6s+T3cv+BnXMgA2gWgv7d0hJl
IQKieaIuyK+bzW4dp5E+daxd3AfBMqMABEPKm5jvxhj5zZ1rsxbJPQAecGBE9jo1GhdD2ljIXyMo
PFv5B5O3V9V9Zs7Tgdk8/Q1kPAUzSQuZol6a/vOWvWIR7BVvKSyBIHD98TYdDedCxnHzXA2rfFDb
3xl1YWC8MZ6HQCG/ES8cqLAAxCT5+V3l7Zuk7RmgAWvihyl87D3SXbkmh6Hvu8bgdmRoQBP/geYW
zPm0zyTpl6Mm3FkXyNFH+vrsWM92ruP4nDHlkCKcYuUawpl1YVLAVDdmLfamQ9vFonAApwwGlg7K
LMsfuYblVFTdezZtSLR6JPc1sMOryvo7CwyX2+wBkpnd1avXne73PevgQiGu7SJbbUErs/xIOMIs
uwjjUm7Goq0cfgyDAxp7xn24XCQO9/7PS+57JQyk+ejlHUbE1NzJaCRyzRbxQJj3uYrX2bSF5yen
wZkPiPG6/b4/ar1j4kvWSQBlUmfgM9Hjbp7zXEP8I1oMB6mQUA0exfGjjouhrA6mDYeITtH7DGyx
zqkPtzZyx+aVC8qoOG+PDlWXkVgKL5pYkpUNC7sbFo3O0vJC0ofva8PF37SFCU6zOpeS1au8qUbx
kadY7LWhorBqbDYBm3QbZHD9Q1DDKqjss+93uqKlgwCeslhvjakWNMNAZeHX0Vpj+a3fOk2L3EGU
F4sMMUUyEkHsBWNukxaKU+eOpitzCu721BGoAeOBcIuzGPNEzWZVCM+77SYwkOousDFQaIqZ3JJk
M3OIvqRg44GrptfLWR5k8oISGcZBNWMdn0U+eO9Z00VNXs8dAAjldVMkJQh0UAye6lw+dMC/ZthX
cw68pgPiKHO60/i6cs8Qv+Jia86IczcrF4jWYV0ALLQ3ytEfj7mxMCAb7FUq/dbEtnGbv0uaYTso
yYa9zx7KjY9YwbFP6WDW26RIeKswdljpBNf5DkLq7Ji1XvnWDYIQ+oaiL3tdv3gEYEP8sMEkqGkt
qPrag5K/8m/2KWpSxq5c2FwtPWKgIMKLe9FUi9EtYagrRjrvlXyQuHCXhXmRFeAsbteKF3Pzar16
ok8n2I9rEc4UFEWVpfUf3K2OHk0EZXILXEH9esaFKj+/B9tmSiVpVwsmc8PTdmqplgKtwKa5LfqP
A43SXwLrXMfyoynAY5KcjTXaURV9C0gHXQsVtYAG6TjO/tPU5jixGqX+iGfVld61QXc0iTLTe5FY
r/NceIKfL4B7k2jgFe/WFpN4t0N4sJW7J0EZoYgQsH4PPCVs8BuaYcBvwCELeviIlzWCUHO8cUMD
kH7OSb3tKUPiFpsf7Go/DOxSCfcno4lltPeFsmxL1O1RznrYXegElIrtYGnmjIYMqJdx3m3OZPmU
+Xqgoc3VXrI2xNfgQihuGSrpYp9DU0ELpC2B61d7PXy0bODHIOsWT0BAXlB/1eSybiDMCudE4uf7
hqD2Tw1CSh51AUcrxOyaGPIpsiN8X9k0ItuvEAMfCKP/SzNgbR38KauXUnM3lxOaVsa0g6k4SIJY
OWBQIwhKmpx7bBroKUodyUh++RqukwBNt7KlDaURLhxeqEKSuwdtscPs2QHtohCratbaDMjH2kEN
dbVzEe9wZtJCEOMd5ww9xozDAVr16nM48ie1kMpVVb4qg1+Fw9GoDrWZI64t7XeiVvlbRytYm/H8
hIBzvc0NKnTgkAhkff7E5kKAjA2ayZptyVltzfwNTNrsp9TfE6167Bx2nRGdZos8wELBy1s6jwV7
CMT0qQXgEw86jk5E6V+J39O2GwloHtf21t8YexQviEFf2tN0PdZ3gEH4jgsCyGcgw1DvVgpoBbJZ
NclmlKiTRzctgILdo9Bn19VqnilyikgBcGabTQ4Lgcnu5kvo8rIVNHWTDYjII2aA56QLu6UlydAL
wPJG0CQ60aJOZlM/rE3uUUrt2n7m2VvyF6MOHD6NpquO6oAb9gLVjUOq+p54OGmAnBOqk0uQgjIT
DfpCwFwETn32pe9HqhcJD1wyMjMg0yMhMJz0DJmQIl+946tD7sQecyjxvxTJ5n0/bKJuH8Y7JkdK
Nv4dzGw1iMZf/9lVfcBR1oG8F6J0U4x5x3Bi4QBppE3r+TulHiP8aOfHS/GuR6htEuoukxYulIv3
JrbJUY5KRqYRA8680UTzU8h715lHsyG/NRQYi45lGOl3Zjg6ftOtFoW1Z5RpPXqw6yIIDvLLsEcv
5nWcoj7WPbICfYbI0syIXkyAJh7KHq8RSx4sJ7eAt1mbk6pNPZ+4nymVXcsToOlEyTQujVbgKDiw
ft3SeHduN+QCyn5Kyg1G7wKJNLA8ZhpjbGy3guZuzFCMGveSnaTfZVzdB4MqrqMPeu+fxEgS8Y1x
V5lJcTFrVGZCe+L4/bQKDI4PnQFAhHZhL9tlanWXyY5hQAEOlJXlCoIUXVxGkqu1RV2ihnjLkmHq
vIGieBZG0a0KVJR8+GnrZsC7RNmUhmqlw5mkNOhSNnLkyfBTG7nRtZHM2sVj6xFwX4/HOxWPKmxU
FlXJt2qkn5jmqOhUxdfx8XBtexsikiuAAkn9BctSoSRjGDqKBcDxDQzm0sMt5qX848CbqjBY76RU
EKFaCOv94RbSVyfZnWC6mqn1A3xpoXFKbpLuhKaWAPurlS7hofzMdJgF+jiDSXb7dQPMKXrmog3K
ySKFPb9490KW0GaG4lkEcN2jfZZS1WmVrp4g/hZ77X/igLMxQ8OLdAXDck6oKzQmpK2sJsGVjO19
ybEtRuf3fOe85Rf+7up270AT8ADviVY0eA5PmojcqDDh7AhfXVrgN/4AHbU0/EnV/ztAQFkRmmS0
NfxHN1EUyvFZM0vzzg5DojgftvcUYt19QGAgMyBWtieUi9fYR8uPMA2QuE/+/Jg0ie5oUhmKSbih
7XbGtACon6WIcHtG2m2WvygyNFJ9twBEiBEysR2BjgHV2NTLKl43uJp9rYx9LyVV4HMpfpCFhhsR
260Jza+S6iOuQBEONzakEbnYWXuzTSz/i46EKKIen4bPam2A+8Y26VKIgHatB6UGkMl+1LO7oVFn
9IfoG0Yx59Ixx4MZ7F5fyPKvvMiqrm0k5aQ/xWIk1Ibtnzt3qVEOFSt1Y4ehA0Z/B91uVoC7PxkK
BAgSSdNteQ9/ZBabgKJz13DzyIVHdXLEY9sXJcK+jOs49ZwSZBEynX0QwJBpyA1avFLRflqTYhdb
G8u0XxNVLLjy9V39JzoY5lgWXjFhMEh9DO9aGvD4QUyaoRaqzcTPQ03nlJ9p4GSX8jJPyfNvek1n
ETXpN/a4rSY7hIvS+CX5n5n1eWvwJ4qbwpusNQcUR8z4FNr5kt9Z8YHDj2qcIlZg03bTPci2/qun
Kj4X/3M4iSt9va9bkHmA5HYstiICoQ1jDS+OlRmi4DCy//Q/cZyqvWmSKr726sPX7sVcXL0H5lQr
5e9Pjv9SgRlGKucKigRsvM8H0qbJqYaDzHYcsyV3wN25RVgBaMDnE5vj+OujRRnlbS7pEfU0qPlc
dAKofmgbwYqg4K+K9e8rYhlPxM0wGr2TCr0GFZ0+cm0GqqERWjSqsbLCF1g2LbMbKPXneRaVCX5a
lu99A98E0gVAWi5N1QiMzDyFhrg2Irt/RopxeKpon2X9qguI6w1lmbEHRjCT3bCRb9GOM9j+gr2j
kUazSlOUJokBCmAv5YtOWZzVt1OwAImG8rAcoxZke1NCQMN851EX/xmEF13gF9Qm+LyXut3U/Gus
ZkwF4GguKU+FnXgiTAiPuVdXNSREPdyt7cszhuZVfj/0eX2jEEAB851e4Qf9Xe4VnraJPLVOK06p
mpyqDNuQRMnNNOsBMtkgRBpkwdw9GyGMuWDcER7d2ylnWWNQ2AuJozSirdPAmNAOA8oJrwDdiXQY
C2x2PJhK84X4Xb1flwg2HHh/zB/h5wP3cszBYqqa1tOV8csOZG5NxH3g7xtC71wvPfmOLz/gFrye
jbK4l0CEIi3V7NAHt9ttVOeWZKjBJSGEWOZiykh+LSfjZn+Js9f0H80IRbg+4CnqjKlpgRmDAJ7h
KMJfuYV0uHEe36ju3dNRlPmfX41LflLXS4GQ1Say/ddKpI9TwyTST3fn9Q5LRkh07/4uIPZwQjln
mZwZldPWFxGbbslLQJ0p4guHxG77QZjlmYLjt5ClY4Z7oHSyEctCAJwfssh+Xh6KuU7+a6fRbYSq
q1xG95PKgif/+QV+xRGjVtKSXuTNjug875xKYp933lSBq54FTPiwUJODqcZqVqOAT6KxrbsVFnNI
QFal4w8HjxXqnwYxEg205NHWr7S+/vWJmJUkfvS6zmTM6te3ve7SoshwhdLLan1kL0WEMnj+KA6U
lWo1iMpgzF3eJYDq9GxllePHInaz9NxvY4ndhhiIuIubHOapG+QgveLIXhAQBAbiRibAwCIJbw8H
1UEBqryBidsNVxaDqCbr3sWyl1iONT4WnN9As8DnPMQlZQjN/7wU3wudh4S/R+rYnnLnHvoDfcnU
mRwDR4l7qVT/npSTCV6ddcryIPBoBl3T+4zfMgximKKFdV5xwpZ+CybvYY3RdMeZe0zwZdy8aG8K
+mPE4BHNzXdmE07TFtKXH2mdPdKgJcOkk05WLvmQcczGhBAUOXcaLc7HPBDNunFU31mUAuMrzM9Y
cjMkbwkhPi7w6nHtJmzPqp1m5kMA3oPp8qnWX9NmtdtoALewyC/gl6ZAOgJO03yPEG8QOhEPnV7n
dhzld2baa+OUSWcVNQsID8V2KkvvhL3KI5q5CgHPqF4mnOGsCumhpr4tvigrf6qMyww5+kG3UjbQ
0p8pi6iHFcP8oZKIc0ziphv1VXKsgTmZ3MXDcmImYp8t/H71XZmJQK6BLSQ3ZbwdJTPZeJh1/LWs
0Tu/vb5U48xBW3evTNQV41MBGlsLk/9PN+fmf2K/EoWaDFfwOnfjfHwz4mp9MLQ2eTqfG+NosICV
HXc4laJwwNXeB53cIem6/eeko3tvs9bIm/gbsYpkeGhqT7YupezdTXIptn8M66rNiAoA0SVs8BjN
BA7cV/WcWpXik1TAM+JRQaNG2XFzAMBmWW9BKDHUShxB2c3zaowgCk+3PN2MAQZ6Jtosj4Sh5Y6q
inYy8Bjc/GPI7KgcVhkrTpc/WVGTCL9uB6cI6PekQk72ueGhbzNYrDrP3AbHDbgPcLzFiMEOCN0q
FrgiBh276UKDN//cdj/tOiDwOs5iROR1p9vAe/gKeT2OPHG1kPYFMbuHLR1mG3/Fv0ko38YcEstc
4ChkwlT3QMf7g8U5eo+PoGkESysYSuxvR7KPjOYeFLNPn7EHz6Xa3thXgZvt2rj70y77ytKpcFyV
aMtDirTpozxscusSbUxdxt9aVjQAFUkcEZ2lt3DCnAEbi5zmZ7LMey1g3x6qtzxURefSzcEgScBl
8uTnyh47ng+vGd4rqyPO1lwnUFLgjc/T7Zv/nvo2oYeoUxH0d7I7s7MjM4LbvjLJ281+YZl38enw
vEnarPMNzAiyPkdJ8evCWZzct4rYPFx8uy/l2ROgl500HNoo9pb1vzeGmUltfwVN175WpSGPFVxj
nfoj3Q7T1RhQkJf6AFXtjuHjK/r64lwlRv5LVLhLTNeyDouOOXai58X0iNSjyIzo2WY4RNwS27jv
VCpeoVbXkYf6GMHUurjtrx9PyHN860VB0dfqX4QlZ0w9KVH5rU+DvBrIJvjpwhUPTDy0Gc3E2iH1
H7Sb82ChC19+N68gkbHFumP7qGx+VuHNZvBiUqcw2/FIak6TmCE5JrM/qOIaotc1yteAPZxe9TvV
eGfNWoXGLA5iCQOi50OV7Rt9kHFIFJemaHbBm+dZyhMr2mKBrtSAyyI0PSzDCLuuD+2WQJr8AeEX
VJ8R808SX3wMQwFMuJlKyqtREWPXqz7aOCaGPnrtwE5wXNvTQpOAygbVPvp0YPeT/Cg6L7dG3Zpi
EVSENUcz0/yDMnHdVVwYrBJVLxH/JfOA+cJaHkEJzjJrCds3awntCpV9ZASFc5GPoYPxTBJz/0k/
I5KROMtn7Rw1wwZjfD9gYUCMX9vrnpyHiUMA7xaXSK7gaL8gXu5fK0UH2aKJkf4yYIlHbkGIIEyY
orLuIBwGWDi9NVd4YOp9xFEUB1Zzh+jdJirUGSKJmijwwfl2F3senWVprqFPoPaIVuRdsY7muZAC
zJotqUSoHYnuNKZK1AwBqYGxnkxHvcR/H38qe0oCCGdRC5XKRVDQ2kUBMw/RZRlFyoVKat5Wf+rz
lx4ERBchc+AsJcqYZV9u2tYmxwmfasJpQ9IZhc6z05nLA8quQ4j1DdEaaC3eaoYwFbGrY/6Cxxhd
tnODXSpZzPCB/RwIWV1eFnSvGeQhr9XhvJn4A4FUHdNu4ALCmNwSI/majbzeHVIOekpdvimZybjd
pmTn0DcQFKaavJwNTCKWqrOfutwFlQZTgzwHHvGFzBlBoxVbvlbeezVYjZ7mymi66/5tqVSPdmwv
UiXSrEsQWNTL3H0B83mRSs/B/1uAOCwO8tZES0LOYSagAZa71bCeMR4jpvCWOJvGjUFi/6q4f8lR
X6Vhi8TOguLd7wknHENmRgIH7eEy/cVEC2FcGOB2Ax6T4Gb1iXQ3cggSERI8EECNpQdUWFMBwTaU
vnP8MnHrryt7AEAmTY2VKkSZ1xk/PTRNrQLDDBokTfblr7fw/nLlQTkRB4B5U/VbSJFqm/O2sckl
l+0hCu5BlXv91MXS+x3bbWRmxCItkYAS2NHfBy7Ty4KKU022b6pMxVCLFIeYe+BXN8InJjxOcY/x
JiqSUDNi/qhWYMu3d79aPJF9jfeK3wF90V2JA5xQv2KK9Y0I4aDav/bnr/nJshb7YMDHD3M+uc0U
rYD23fC0HrYew1mQrOP/q6Ro58WgIN1PbmSWcW9rwj2TwjKMHRB7KqZCMso8WYvok3KGZDkyl8eQ
6260tgzLIYdQXp5iatAKVB/WtD3u2l2EIYMQzMAQSO7Ezl0SdPnplzM/+9FUtu6thFRZzoS+uLLX
z5k7LRa1oLwXCeqyvVXoUJXIaHMVeXe8qXuoMmDJn9+p8fVP+E1Rrdtqu9oNZjdqsPSQ+vx/QV3W
f90Sks2Wf2JhBtzzfKNk/XE1ZSHC41PA8LTmzb5QwxAkLyUZtkLzJdPabdi5CdMDaNg1qBkBXi0M
fmSxST0PqXTQxe1E6tI/q5HTDUE3Xmp2OhI6YpWrG5ZT7mAmOGgkUBNKfQX+XxVY/Obt5fTA3MmE
wys3j9PF/2YrvqVWt/0WO+uZOM3aR6rdBDlRVP1TY6Syi+MNYvcLm/MipG6t726UUCitr1r29/1R
gqrcertuDn+QjP7epF6kMvjHHqTtJHR5eqEroOYK9wIuylgQM+zBgo+r9UWkjyEfAlndtfEX726g
6KcJ8YgFw8c08IoO71nfdnv9A9EPnIobkeUn8X/ZNCwq9lqMmHvGud4X8D0OX7V9ZnzqmD4JrR1+
VWiieHO5lSYnFYLOjjU6w1snDJY9ZSNLXMozQIomSQ328+sPaXAArNsbtE614QzZv6Aj4gyNmYjc
UBWhjATO6ipHi4IvumJoytKzzqtgN9AEA98SpTt1xpLt0WjEt6yN2XgRT5zBUB8GgoQT7jCyLr/2
7X3elwg+Y3N8X3UVE6re4IZKhjenCje1OaiJbEEs8iCzTX/x77Drm0me1NOFYHBaMfF3mkoZ5D4b
BRak2Igy2dNHmZ2kxOKLFglV1yvhTjmDuktrOl1Zadyuxh9M1sKEmSSb+Vpo1TE8VSTn6SiQX4yh
qXDG2NSar69YYrdMNqHC9hlMS/k/NaDaieKTuoZnTZBHdvZvC8nCHVPzFr+CXRkZZUcxoZ/WloJB
Wudj47glesqljcGksVDJhvaFzLfsEI04yYTjhMq2E78oLq5ikdlEOirRsPTiPrxI2+GiVWw94Ew/
a+arxGbjfhq+VDit8Ol5sskgdVHngDTInyxGL1zWgRsQsThkK/QbjJtRf8bCBYoo2s1rmT9TOAOD
mgftDI4jZxIH0EuOGjw4EaUV81sqqiGfu4qVJzsQx09pJ2S/wmMwfrvIYnuq5U8f2ZFxJqxqv7q2
TmIhU0LKWf3KKuudvrYocWMDp09XJo0TVGp8nYKTSBESqyOXpxYXhouK6KQvMb2zu3MLpsJHpC38
4XswTHFeBTTtNjKMV381jMn2eoKR3kaSOeT1ITAS++ICBId4njNjM2Jy/f4QSyG3LvuL66TOp27v
hHIN7lHAPAACYHCKWv2ThKO0JH78Rvp4Dsb9p/khGDz09nu4BuQUcdd5T9ImbtyMzZae1ukPCQzi
/IGCsXI4MXEhuVFGFcwKiCHVjeORtHveAIqUB05EO6cGcL7FZrzMx+yXl9khCrzYBs+vxB2hlgrV
ZDSr/g+TYwSe1d0ZjewHSnZ/HV9Qqhxf8ZcDehbigYkpxsTcpZBjKiEi/0vNsQxMoP1ZWx/0s0HO
wFybjgA8iIXrc8mpqUtbfe+KVdIiUndPLYaQPMRFwJJx3qf844hAIgD9Tsgftfuk7yr9F/nQRD6l
9BgKyF2YzIAoZR//bD6EOZ3+OuFpgHGMjXJ0BCznmTkjx1GssQoD2dZYlKZmdvJVnRk6xvFGNI0Z
EEQ3ebPdMgGA9ww3T1JBBt2pgnBNx84m90b/zkUtVBj3BsWzpvXLAXoIDltVD1EXmTPgTQpLihfs
k9k2H9MzmxqQe8EJkYkiwIS0cvpufchp6YoXtV+F4CfLtzuA47s0qeTFCdFOehusyBl6en4Hqp8d
9Y/+2ivnzT5c1gx0lP086VtGpIinygCMCtci52/EQKKwJZYaDmW+mTpIBhRFcmOLcDI6cwHa4fMH
FUniO1UYwLpsK789H7/MAmzPG+L6WyTTVd3tPMmZcEyPIJS1g4N+fYvXiVuhJ3mbDSasrBRvX+AL
5LxcjJTELNOYabBZIjzj3wfvhNvWqhgOPbRJPaELmR+OBsCOD3O/cXnstJWojO6mS5iUJHsau59g
ZwqdrrnClXGP3vDKwzxQBft7plVZ0yg9Vx/Ii6kNvyFfELtns7MgUzE6dIIoeYhwDLwiEvCeiTgH
VXzYVZ/goYIf11IxtHelfxfWMkGmFvkZNHv9+lzwxcanYQUXDWNHEr1zq2McBbC4grnZife/5/ko
mJqMNnrGeOKpbHZe2x20l5VHvLhwkAI0Sc4YJIWnowIwYwJVz5ItRzL9Ard8NqQvrKbEIiIbrkbv
Yjxp6eOzKhiBJwIt2TIAiGVgeIz1Ni8TwvSEBneL3wpa1l5NI3MtmIDMwvnb6PqVRWHHn07yJxrm
KgbbbAP9GNCTvbJEDeHutMWciZwNnruGgnTYbqqf/nAdMKVgfoy30dKgRdmhmiBocP2ZjoHG+WdL
Y97WxclE+3/SsOd5Lv7/RbFQBmwJly9Ls7XmjKWWj+Dy7jvtfDGFjC5jn9nHzULmBfJfTt5MvvQ6
xaIvigUMN5FUHQtmzzqao2BzJurZuJJtn2HOUvtF5748FIvv5Nee6TilsEjJxOrsDRuqRI6ajQmt
CQPyEB8b7qtGXY4ea4yga+ScEdkvor9E7K4QBTgSvIryVwMA/MgJoUtBfumpWtyBQWJLTtPipvY0
UH/3fxF0IJhfeeBYegW/v5Jey7OcXTpyDL24VyZoCOgji89wYE/ZAiQv6HvCSlGdn1gwZlsllryk
MyPIsV6tslnArU8sGs4VQkhvmeHu5js6IiYSaBsZOQMTV1aTjDp/WFFTu2UQTkCa06/lpHnq2K83
nC2sq0kSx7PhVWHNUA18Wo9h5y7TV1FQp9p1033r9yNr4WLcMU7LM1GzWa3LyQ/mLlqPrrCXkBDV
Qz267WiQfqCcyMdd0j1CMQEWOeJhgXem8NcKcOMCWWeM9ld0V6dRZnwV1MCEx2sM+5NSvhojB4iK
DH0NFJP6ZNTVWTNuqJEt9yJjvmEOOfbRAny2F54mu4I0iTBMbr0xkVyo3sxQn0HKo9Ef68dO5Vtd
m7NbGdcJMzMfBHbmHqbisjyF4a0k8sCGcVxqYdUXkAm85Pt40/MgNVnsabl+5cvl4rkOY29U/8dL
1wpwvYnl9JU39wQEuh3sfj5p+/8b4v276kDzEZVfPD7593GcW85tsbnavvCU5D5jZGZ0P1HSo9kU
Asor7rncftUfbl5/0yEMTZk321+8yw2BUP2AyDD7Ak0WA83SbrXQCpIwp7iVCEA674pjFuo4SrY3
n/bvCz9f9lPuIn8O8FtC2YvRfsJbv0lQRkLUnHAsxNIH6/nR27dzvrNv03QxAGiOo1aqUmXMf+J+
YwPLJi+icAw8xNY2c9gCEzRRMi6uzeoPrzKFpxSfT/O9vEp1DcfFJxMC34YveIAuXYqpGUIRuKxz
U73QlxqJVtQWlt8mcNAIrvbKUgW3hdLGAIldqcbksW/IooE9TaL38qlQh9m7iSRfM0O7KaiKDnxY
2PQ5IejPqT4vGvHLxhbYdSKPsu/iOJW2uzoqcf1MbKrH0hpxGmHOeqMJ4mnLoMYpdH4QqXWeCJBx
57aTNUlHQI+9DwxUuL3wPzThp7aKsizXJ68CoPnYZnguN9cUHlv2gbZk0gs33DlwrTC15da9jy8i
OGOOWWmNBmpnKYY9C2eJPOHWm9GphNsfeiFhygUv+L1lWiWvgT1veRzvOmpFV0Vg88TazaDsP85w
YEEX6wx0BHLNLJOwKnc6Zl4ZGsern3mujtArXlxwQkJwvshf2eRGN1T8w1fW9YGNxXI3rZj4qPeJ
3luZBp3DDnho7om2reG85MYXLQaj+fuxFScCP/OUkiPpTUnwGberCnBoes6v4sHjyph2AcyCLw1m
TPVEjJbaXVTPnTevulQsSNBScIA7hSNIb3guqqT6CJKz+2mrwKl1UoIE0n9ejQKny9flFHvA+NjC
Jd+TuEJKQX4BsOX9sWHIBKO0Yg/KiYjQyBrjj8lf/HerjKwqvJt+ukY4DZ0iUeq41Jl5FiA+lkG2
62ptiH3avknt5oQUbEqP+Q7okmAWc3Ok3MYeY9YAF4rfwduc32H9veWmIbOrJVFkjiW4tAcvN1WG
/+GARuH6feEH8JpcsWUeHSz4A6fJ+4UXl94KKnfMZ4nppql0O2M4iuGrSdHJUATqIf4iP/xR0acd
4Xubnk/wuSCB82nvKHrRldiPYd0DNghUUCXXbnu2Yn3MLmYcb6m0thBZiYRARtFqBM+a+CdYyEnb
7Ul/kAW+7TW4trTN2PbsnxiF1dVcpwqgxpurmhHhNB8maN7A2v9UI2Bh+Ek0nJ7tITKCIhtGkEvZ
1ucrUTLwnyTJac8BczPq+Zre8QiGnjlVjHBY1mnJabUIIG8TBJwfwQ4EeliyXnkDPEPRXudsDGjR
HvX/ctpYHERAn9yzQe3oQwBL1xuVBrz75Uqegb5nAcuBcMDStFxSb/YZzRw6lYeLd2CxfKJ4kYZB
kg4DIiWsrLuv1vZHY4GGNiasPFsXB7YpO1LA3w2o13wiOsKoPrNaqUX0rC+NA/YizP8zw3IJCrNz
xA0h/7CI8kEdLKj4RXTKsSySEKhICSK9skPPgq331RAkC2Bhjn7SB3RhsGysS7ehvAA+2QSh2nnP
0JomzX3kNzXT9Mr43KhvhjKj4gs+UajrMJY+ykwfRZanLFYUmRHCJiCs2Kl1k7u1UMyatAATBKlo
B51w+xSGIgjUOoFqBD+KztUIDqJ++Isd8PXSFCiBIKv+WnSycJOlFKWmDAoKku8Lg3aOBpyVHtEW
KQnsUeJp/U4K7nCR/tgLuB9Gjm2z0iABRNe5PAEQH9HITCQOTGFlqa+5HvXYkGAgu7BXQN+0DOAL
F4LwL1PSBa26F3oGHwbP0zQTjgJFgYO6eMHz2JwHiH3CAMMll8JzJCqSENFDoWdZk7d/K0s1+uAC
QojTRVzLweOsNnMRx/es/zV8SWd3zRggXmVNSaGYfFgB6HEDOhQ+o7rplx8d3Ti5QppsMRsrLsKD
S5opKCp01CCJZhuC1VFq0hf4ZTyo8A8QpQZNW72HhBD5v6UpZoGGJ9kJx3tzigWBjuzUwGbKa+32
s0A7NBvc7ZA+YY8GOijsG8lEVJf3og0DyjTIWGk8d98GgYWRullysYsg3fIn8SnGUtyGAAAISeFO
A/omPRfL0CUGawTLX8oE20UyRCGFp2aXyIvBTexJ9eIvavTHxDiLnpkvOMyozxNS3KkMkRz/4hdp
nwctMOhavwUKiK3NbqKHYs+BfPDBflCgMjmtzDt3hDdkqN+KEW6t90G7e1DOE6yrIoe7+KS6yKEo
YjO1t3mPMJylyZZhTqHsxXFUrePOyGBORBTydlRo3dQywQM8qXCTGeLhXR78xkn+bVmsHkITJwIv
1BeWXfyUhxIUhF1s9YCC0kZRVGSbykmAncZdHntmJFq/m91rak7okrV3qelV5OirQeJd/SXTzv8M
Hel+gvwBGrEVLzRCHbDhpDk5QBlz/6dVgcE5zKCMibUn1Ryochm5oSkSFyOsqKR5TRxMruMEW3eO
w1iXB8bb8qhRfl2AkYDcWGnHF0Lr+z1ciyUyPpF5kj186HBL9XvmWxkrOuDvWJ6Opce0PoZKOacb
4qQeZPRetMOx/hiTGPFn3+qI99vcL+ZuSpVMEnT16UjsBH3ouFF3XANQSjnEHsuHvmk8qEUhTSOZ
yIbRUhY1OikMuUFx64Srz8+NF9YJCCPo+/sKt/vxNPbTg9i6TKvuSJAdzcX+xghxV8qaQXLdXxdg
l4CqRCaOt7ka7zrTf5y4LimVVi73fUP4VyVLWgxs8ci5mQw83V/evGxYSK1hwCf0D0+kW+uP8cKR
Mq2V6LspiCQXTgh5ivqDnE5wIC7pALJv0VbRBsR9JxPAiUKBxJ1kIKPISINg6RcYTsafmg2VF6pc
FtbFR+MyCq/RHiBM8hJuf7/OIn0xl1AVGhbybqcPKIHCaqk94H6m2RbtzbFz6CUfAsPP4F9dziqF
dtQLpllPUzLL2XwhiR8QssZDGg6KMyCxl9jSR43eFY8awz8d7jsoNutJuZgVt8rSSZqqtrKzC7Tg
2GlYp3GFY7o7cjxBeL8AF1P5P3yNI7KN8lP1zmEaAhMAeQVpAHDsoTOqQf/LbHlOfg8tQDmgfsSr
OPTsN99ZwmIvl4t+1v2OKosOa6qVNgNa7Tg3Wq3gi8SZ1rq4oSx0EkE1ilqG4oV8zU5wi3Yr4rVH
uTPxHBUjPMDAijbNgVb1VylBpFT0dcY5UIAPxghkD9sImC08ARPgBklIGcJarSe3bz2O5gV5Ri/P
ZKw4sIT+xp5DYN30p3hZSdSoPBsQkVeVAUZ93WfGFxCAI/lNecm9qTZl0RJdZR6oBdo162/Z6vNq
WmaQYfCW5jhYpfxln9YzrGJivJYcUCW8BIa/B79MzJPsHQJaz8qrPnf8Vur9AGVctyw+fx1IeX2x
8PNFIJttRJYIQDcfj7asLq2yvzDQk4MCIfcdlIz/kqUOJIY7Kc8u/+YVPpTQkkiQE4R8dLcUEqg+
QPB7tjGnSfjLZ6QDgawXHxs885TGEYtoBW90tFnMgsEJux77OY0lsbS/K0zPdcA6xi3wodQLaqUc
PTFUvBTKps1rUJvC8HX/kDck/iHaLSXbHR3Cf3zsylBZqthPafSPJGvsPc6QGI52lVeEdoTyoZC0
z6D76Vxa2mLhZSmRSUJWNSYTukXxIlkyWpEhKoenH4cQFsFOmMyTLTmyin2frkSY/zs6Tv+RarIH
VVBhTyBVxwvFo1xJrWHBBXeDni0T8HnhgwgzGpCChzy7ayF0DTRtlhWLMj/EFb0sMsVaM3UVZBB5
lfoF0lfacL5bMDroquJdJglU47EnTyAubY/K+7ylzisgVFfP8AmAGwsO2RPWnxwaWN0nGerQvCMZ
65IUbaMW5WGCXvOTxIg6NwZQB7q+RqYuHkytT8JCOHcfdEfjd4Juv7bd0PKcyXjNu/9x69HylM2/
YPsqRExHHFHVTnoeW1Yb9p3+4j2X+PMFblLTkHqRisEQt8+Um4cwULHh3XUdjHnIMa05g6l8pGtG
X6et8TEHl8SmLv1iUvJ3/S38wmPupy0rVuQDMBE9Y5vyrFB6YwsDF+olin6vsB10X4fQU9FN5v2I
rRyIroThFZxV9NuZ4s2kLCRkbQPrX9AoJrtUJDstXR1Y1ca72fVa8DsbmVToEvY0tTfViKbuLCk6
s60L3+eXwAgzxdlcnIu/J72sYv926nt5FP02HvtqkyVNaphlHrfti4GMCHxtmLFqL7g5+kms8Sef
Au4FCSPjAn20RQVaLPrhGk0dpoAwKWuNq/+JKAWwjiV1Q82AQP6uO0TQqvcGoCUTsxHqYESJAokC
Pv/k2c8VHSttoR2AYTys3yg/31A9oV+7jnjkuT5T3Rx3b2J33tXO1Mi0j7DJYXduqhdP1MJnneln
oZ/uiznbrMto6KjcxJXZlyfijrj2CqKQaQIl7mFoc6JD/mJHkL55DClHH03YkdM0E29IsjKzivUL
qN/C+EmGmZtCpS7MmXq8pO2P+XBDP3w9rqTNJoEtB6ZzLcVAJaXxjcm+HR7hCWPEHsn4XtKQupFe
8/vmRzoN3dPJpqR0BbM15mGgI2TkfgYRJRRL2ewuvKgkuhKqXYcAtwmvEf0DJA+y6EwgFwLHirLN
btINkMDrWdSD/Upe76BIt9dFOP/u03545KE5yVGa7qCG3iQ185i93ABAzONrI1LueUXuOYVPhY1q
p2sCLloD+tKN3ZZWyxEE8qVs/AWr/XEJVnbBvOQKkMRVcAwfr5dV9F0T3nSggoiMML+sSVLTzgMt
SazYuxLAIhXtb+Rj+QqOky/JIgmX3jpaHYzTHPn2CXU0NViqAuZr5ikrrxjn9InGo3TQsOmsAKJ7
4AH7kNJl/JwUaSrBlZWuOGnOSG4Vyd0uvHaFYY7oG3o8eQpvLScn6cJJnBn2kIcgsVeoT403s5Z0
aij7vCxVpaFqv0pIlehW1xWgqW7TQu9kTPC7d+kmkZ0OxONubKRP/qXHW53Yuiiymve4fIUjDlsJ
xOk196Ev1HTGCXjxT+caYD4o2fMCfNRPhv6P/0Ookr8W3vdLYzr0ENuymxt1DZgE1zrVElV9k6D4
RfoqlPBGFCOj0XZ+cbm1F07oxsh2AFh4I/SQrLE/AujVCFN81ZeFlXH1QzWv/xqLrgngaTDCo4eg
RbqjECag4n33YOAfCRRQMFIZLwF9dGptBYyatGaZ+gDuEf1h0szxC9r6j9a9Jcw4rEEVw2KFjdVB
j+QQ1Oq4n/isfIoBBM/FEklY/lIZ7gB+oD5Zx4WNg3unIgGHQfqn3G1oXHs4YGesoBtf4W4eMM1x
m+QL7WWIQ9LPkMpxsUibTsj5VWjn+r8Cv3mFhet3Gk7lW/uS03gxjmjNB2W7wtC6V9UddQCginta
E+8jXPiAJjwhNSEL6jtxkLJDescOnSH8bI1o+M2fekLg62O3hOZ9emxwv430lDxRpi6wlwHRAfFz
SrD5EkfJmz2gksqBhv3jacL6PddpcXRHD67NF8Rjq1Hc//YEBK/i7qBKlSy1+EZ4Eh5QDO9R1frJ
tI5+nxrBSueJQldAnyncB+hdrDNAV9hCb6MV2saLEKdR0ZdmZ8sAvwt5FsoRyLIB4XTfO8mV06j4
bXAoLfgVv7qnRlMWPLBBgfIvZmwTRm2J0wxUxXlzdkZcx+FMTAtQoAssVfI3Rthtr7dgQ0HUhPvw
rVf2clx+9cSPrbDVyjGnUtpGUiDtd9IJOfVeNFWlOQWyTWmwgo9mXpF0654t3JbQHfOZTPi4i6Q2
WmbVbdWUgGwAiabdFk0JC5v0Eg6yR+ZS9UyZHYAgoE+jhWAMWu/aYvLa9CbUMCqSNVpyeBVnS3mu
rMBQP+0nSuHPrJ2Nn0FveSuADUf0ueXYJoCuUr/7bvAIBjRLyL7zvYMXSkyKA6ZUT94j3Gwfs8LS
fVKKUu22k+9WPk952Zyhc0G1+aVKbqqfiQGmmpuOFGMbNpf2C/EwdsnD6jwenxOS4ryl4a9SAemW
nFVpMQgGfngWbimIZ1sATCf/BqLO1yRwvB+zKxvAY/7ujaShO/CnoUCpQlQutqrC4TOmOnhD/M0U
+ziPHoxhqenbfUjstG5kA5LTFTW4Xm3Gg+qKbhRPevHCvqY3ZKCcYf2BgdR2OrJ9c4/fylSanqqK
Xxo4qFXaw8ZSl4Gd+Xfv/gdL8LNirv/BOxgZvnMqs/JAyS1BQ7fdIiUbOmzWYd9lMYkSXIfq3Nb2
T/+RcDjd7+3V9b/AC4rG28y4Hi3AeTfc3UXs/F1t85dU5XWo6uhfM/7YUmRdjzBC1vRZgsfVsyF6
wzYlxQHgbu9Ir3IDKiHzJ35NUeKG04WyiD87/bE5EzX9XuowdYDF8fo3mBlg3ds451n9/TEp1L6i
D8HKq9QWnpfAkdgc8tF7/uXVNQZT+dHF2RVimR/urlSJWO7ZXBR6WzxIPnTpWihr8DLZzr9XIUuH
Sazjry+7vpHnO9FNWKg2Q6+ToJ8toFNBTaT1Vko4lhXBJeGJ17zlucK7doOoG+Nscs23XGyHATDE
qLKCvFZDiGtBS7IpcJAuXCR/71j9CcJP3YgBVPaW4sFuRLwM0l1ImzgWOw8a5L0Xwn0k2fmfs9TE
pdcI81AyUzomUfnOYx5w+1CvIoMf5IEZPbzx3pL1XjivVFK7wRIRkhNDGg54go+qYWCu79y0UhLa
3LAO1SMGOhHU49oLV0+AqHzdg/BVh/6erv8G9EGG1meE2t8Tys63CzdN5keWwFDHp6wWZ5dp7o1a
eI232unyU+FLPn0v+HBiJyl/543/NqybagtU9sBThf6u7qwmyX5CTAwQmdv2RRMn1SzoAaG8jVvO
7gPLZcPDhb9ePDeH6HQGbLShV78YOTsfhLAxuVBFQC34hnfIvz7ks6vJA5H8s1tC0adHlBdCtMIj
aIXqlSQq0UqFOEu1rQXnBGHdBAg9wzCEL/Jg63BoC1oTsryvivpWj5oukQzUStxscBZxado6jIwY
gNXpqL1K/nVHK+8l+nRtNCT9X04fHG3IOHzMgx9yXz8ZEaaLcdjxz2p+e2inkCxbgpRLcQERkVry
SVTj0Crx2wmfn7UKnsMMe/OoAvPIBxxXR2F/kp/yRPC6m23Ii0uvXSsMNSRgjaGxLv6gb8GJX5Kz
XrWj+JsUIUgppqwUU90GeIFdLrw97UJfYL19O4ALoUzSPN7HRiObpTFdanhVFSkBjkdcQXXI5Rpa
9eYQAlbhA++TRqBmW+u8W6llvP5BNgqrUfg4k0BZFQ8ufKopkoOEINxOHX0WoOc7Ctrj+N7MfYR2
KEt6wo46w1u7vei+a8TR6Wr3w4VVJDZnIbw3YTHEzy3tf1NF4sh+IEE25YyN610YeEHes7jodBFO
lmdfvQqlXRLjKPb4HdydJdT1T7UQNe4xLZncAyJV7qto1YBWMj5dbYcXGOpTUJB/ravfLNdDQCCf
Pxk327AhdIMoj/y+s/hYr1sSQUY1F1q3DhEZAVDYnNODKFkm1se0vewrcr3YQ6pyebOPjhYa6K5i
wXNswq3N6WzV0LfziiPz5VnW1URKRZdelnPIlvgCeY9orrwbl8+5ZofHoQrRTXB2puFJ3U3Nd8cC
IEAhH/Wjc03FfRjadZEH0GUnE2o6St40qMxTXJIU13Ta2TGdltYwtrhZi/6eumja5kAqLDQ4LjaZ
QOmFjXRD/IE+PEv0L4FZXvh+n1AL6b/gAtV7UldvinlFTwQCKHL9o2le7u/dFZfP6QRNcxzrlEFU
s+ma3jl7+RGTXhMfpW6w4TTn/Tjyg2Akfp3Mbu840A2BOdhLbb8mmExL4AXd8FePpPENUR70G8dO
bTG9xiv9/h3cnWltDCsJawQOCF2ZZ4Ec0xX2KqCml3qWJZlCDEQwTD1w6bdu2CduwqBh686SC3Af
OTEoz/Vx1kMcV3JvNASXihGrQPVQqgA+5oCFIfuHnFd0/sjxNh07r0vnm53XDLO9owjvV71UyxcE
aljbu/nm18I+QZD8n3PAacyIzZz/M0PJW6rU2WqAYKQgFQlGGN3ObN+6/Voh7YIakQBweztwSPSu
lbZwnkbZeWLai+UR8TGwdi1KVPfq7JBh3ETwBdjJPeIBSv19FpKQSDmt1rA8JSgqsY73C+VTUHg7
7UMaTofz0PjhpuZZ15rTpBnxp0LxY+GNbzij7NLMdtu2lONt8exFI1daAwuOpi2F5oV84Rs3EyL/
xs/dO1AI4g1znpatlekMjwmW1Gn1KjNQwoW2MoSkqm02cml0bboF55bW/E+TmV6CpwhS/1Qy1Wr2
ScpC8MUpVghQu+6oY2nScU96a3+fOSAd2UdwyazJTFcoX2IqKJtH3i6Jmx3QlAEKAJbwHv3NxJ8k
sBHF2irA6vcbEHVuDMA12Di83DTUUtHC8Gyt7MxuY+l05gU9+72J6Jh/QJuqEi81ffTE+/btpPyd
zB+gdIAFWtukkMn/49UTru6sm3X4OQHB8DfmBJ3ioi7ZhZsa+LuQRa24xE5Nea4LU4SUL3Wvpteg
ueib1CmSXUHt5AAithaWxswgFmSdNEvxaO5tNWnmEblGs34/IZC6fFaj8gO8rWnv9WR1smDhAHPY
zKq1QBw1L/7EQ26932gCSrpJvi7eNJQkpJ+eLAaBpoYUH5Txd0Uy+YWk60MK2vA8lVAOl3C6akNd
Yaotlq03jlMZiFhpufwcI3RSlGkEQQ/BfJytm+OeFQlAkHKXX3HCyQ3bNp/B9pP7kqG5xo96Cr4T
TeGFNz+/Lf01ia3u+2eBsbHyzYchPKKpGzl0+RFgj3hxSeVAW9UvReA6PTi5yp2O0eSL15YbZSS/
0O/fUbNlnuZ531psUsw5ULPk4vA3db97IXYeqF3TMjCnDRG87TUmQr0OODuQuUIbYc9RM/t9JzM6
Y9Ox0AO3KiRL0So6JVyj3BIMEvnnXAcvCAtTEYia8ahSVPvXdyjpg/J/uVS6N7fc0yZYcmnHtEGJ
cxFFTJY2qoqNiUSaejUeE9thJuuW8Yw2y2CpgcjMo1ZYK2NdJ+LUh1/EG0v6sgTQQxgK8qkomu8C
/uTvtF2bVskqUAA0Pfnou+SBPmJpkHlwC280h8RV3B4zg/bNGis0tgYFAifvQ7BysRMVw1yhghdo
Zews6CNzIdGHBYetmkDknwQaDHSAVQrf7/aQHrkhgjKq21JSF9yQgnPqdMYY8oSSFbHpIGdrlt0p
da5uIiB5kcEHzBfoBZpoEh5wmZAcIjxr7DhfCsD+NpuRoY6YAkCCvrgThU2JSOORSe3JWOwl4o6j
kf4ir7SmQ8zI36kf+qJwgmu4SsGjMLRU2W61ncOHLGK3rGP5/52ZmFTthptfTInjdPGd72HBq3kJ
ljHQSyzDWPlPm956E5COb0R2SZEGG4YiyQgmu+ZzNNaC/8BkBeX0I/4JlEjyYrdPCH7qgLXzxbSZ
JOmaqtCGLA9WaVAG4gVFs4CdOlMXRpJKtRqCEnPy9Vj/wMAAp7utf2U8tVt2BDxKseFBzJUCM0rz
dE7+otb23SVzxtmZKw1xd5dttW6/BC0pvSSUEYOUoFi1GPX/l1DA6gPUwLmZX8Kz5fdTJfVOuFuK
e8T+7DQsUaDmeVCx6RNJQ1SredM83Gog3hDf9f4St4t93zOC9HJKfil8VdqSOwPUyc9xhvT9jk9v
7sehcK8ummB/JwlIdfdfy+J9Ox79efT4rxBbyX3sXbvUqZOu3sxHj9EWRpqYGqxFrDL+ka3/etPd
3io2EH0O/U/D+QyZ2YK6QetKlAG52Pd61cwUKYxQ1cKQj7dTeEa+rWh7re7nl6lbmHtxrh6iXT6k
+kOxcEtXcOjV78AZ2nsnCZC5tkcQ04ozBu5ZfCs5OZ+fS9JLeiKduMGDGSgtUC7p8uhoMNORqcFz
NFE+GPCQqotOWM45BBm9+IshEUULJ96fYKdakhC/BKtODJIzczx//9gKd+ZYnHeqGE6IJPOE/i9t
U/AM+Yk9YIMACjklkqU08QxJZSyd0XLBRO9+9v0IPbL/PrRRckdrxdet61BTHhNlFQH/eFHyetGX
qqLdRwBrpJULsfbt1Ktx3vuFd6pz8OVgromPfM+swsibagFjawEMHyR4TG/7i+nch9t+Ypk3KGoQ
prw1FllvSZT4QoQ2ZAc/YHsJHcaAsaOaA3JEMkuz8Gys3733RZF6KLa4wR2BKhnZATV1VgGOdOuZ
fudAHNL2OZa+OY5OSpL252tWRCB2Vsyh9IcGYgGyyA2DYmN/tbR90Ahmz63dL4B3pfVfNK6/RRjj
gGeDW6LqcmzS69le6kyWld+dhFvNy/skvflpM98OpfaDhuF6XC0GPH5RayySza2Zm2ilUxroJTru
csw8cLCPictVruvHbgYSv1ZWOHytaE55FAQUhh3R81kgiirjaQfwrMLQWUkFVExUV37NCAvDtUZE
nMzhxNHiDKrPPQ7aRQ9/vk9xQkz/ckdPxx+JvY0jfqnOhc7Fts2AR4ZFsE4Z49jvr8dFiljpmQkh
msfD5wFprjtozptV42oT/iY3pbWDCDdVP14iMnbFAG/OFKT7MmQhsWjApfNa0W7lLAQvgqedRMtd
QABwkximlBVq6Nfw3m4AbxWih0Vgx85zXEh6RcX1x6D6yBVdldvRhenCMmejxirA+bvBO6f/s+ol
esDAhIB7/KpEFRYEWIDzYGH+Q0YLnLVfvBt5L9BkXY5yKZUeQdY08XgNVLVC3Fmo1XCCH1XosunR
FFUAdsUVfA0VCh5a/dmSE+68RhEGld9flqEHe9xxxoxaFw4f2P52OITBl/VKkuclisrGXEzLH8oX
uY05TTg+ZfncOFvo131d4lZmzaxijZy/RKxh6wLHosc1KtFquC5MNKNNlqXz6XPg9zYstblhokQ2
HyV453+QLBztgomb4NBvoenS3TBhiNWL/yZIiG1MiY46CmipL9z5zKHgIpjgeKgf8mL67P42hYvH
+rZP0Gx+ayKW/d1JxGQM04Gb+4BY0GrO7Px4cncbaMLqGBaJR33dAYbL3x3u6iZv25Q16Fec+UQd
deoel7gsmSpRwu8t+QijyAR+bePoUqZ/11DQfJPZ2CVfKD46x4iuBpEPJ0tcVcIMhheoIW2gdAka
Gb0IJDHrDN4cY34PRIpbxEOGyiw+F5RFATiYP8tE6DUdGOKhpgqOJ5pmNOXqxioadtzMTl1et5zU
XCPq9FrM4cslV1JmBME1gU6dwFN0SOI9Cu8K54RMmQK1Wb5N0qwCrLsHvZIk5wa3VoaVYmohSgdC
SQ8Of6lc9CCfOFeRWs1f/YGofzyaoCiRaG0H4/sSFOsAkT1/ECqYtfuvJKZaly02Cb8fo/hH5pKE
5vhK/Z6yYFFFhXJqfLu6AO+OOA/NvGcdqejRDEfvG7t6kqu6kZu9cc1dlnfxJW6ozOCk+cb4htsX
C5eiHhXJWawmPmIn94pmxT4I82bw4bbq5yAjUOJkIRUZ+Nbh6VqmFz+0vx6pBCo/7rUpWDJd53dr
WXLn7G4q/T2qsig33eKU81vAkC4iyiR98fi95haWPKQfO//8zAtR2Aq5x783mZ5AgAzn+Q+gp4yi
triDaQzQo+oDOtgi4q5W8TaEBAVNvjUm8EWSIOSU4ZyA0OJ5ogZnnwFwdL6/EGMJHyud0WJ2Ei0Z
xiQ6VOpTpThHrUNLMRWqz/XOPORu+sXlcsMIt6edOGILgSbLg8X14hgA9HDwLyKZGhAEJWLH73sg
f9BrjP7VuG3kJ6xsijqNEH9aywtKlmFeHARofpxxKKhGKA4uU04Zfv7qItWwkNPP5+JOCrwxG0k2
p5lnZ1V7wUb/rAzs9ge2CNRLCX/rHILqbe8nxPEyKtn/xTPRCdxIUwqv+t2HCOeC8U9cRHt8Z9jv
7owwHYGMsZwdG53BeYPBk3hdSa7Jz4j7XMx3TOKIVZMoSqa/hd5Q3UGWTpPs+J8D53Zww29bkz5M
sd4uOVPNMg2kYQZIy7nZQlYA69Liw6te8R77ugt9mz8R3WkxqAd7U0xhBRwJaIZLMNW4KdSiyJXe
XVqjDdZQG/RejZVmpzUD6x+icdSyjyPsArJkLBiYFzu5ISLZpZOoyL32Goh661kh4lMADpiZ8J2D
JCcZ2ipb08nuBer3Je55CfJhwx2SNUydFA/f9UztKMt0LikhTc7D54cK18AiZ35HigpywDvE86ty
9nwf6ffANl5mZ7SIWWjCmI1DtiSYdyBZ73qDH5s2o8HPIpfqRqwR43FGFJNB9JVETOWcTdhqZhNg
44MulXpgpsiNiDU9dCxWQ0GLwTWJPxOdpxnetww3sVQzT8VyD8d9vuhP9iwRLZqwYtuQ+tMnqTtn
RBVZUu2ayThxmh7VcLxm9s/wFdGeQpyE0Op3FHyLprLWhEjyCq0RajaWbDEDX97RIrNJQKkgei54
XSLVna8spPRfYmDFXtFJHpO261F8nTcKme3SGkElXR6g/fCM4yuEr0EE+XHx0MfwQH7GqdyunTL/
lpVTB36U/PBuvDpinLeRDIEinP7k4WELR/utc/E3QNyzn7Jdf5/YDARCBZ29u9NJmrlrQKHQgUBG
GhbOJGArOcxRGd18SMUKcJsRmhnS23o4EO392fF3bGh2O5TYSiiFUGRmIXjddWCNCmd75tRQJ2h1
Dmnv32phOsZNYr7U5HEL8IiwJQxgd9D7QwKQUmc5SOm85QTEUUyyHGv73tEu+DoetCGPwvyxMyBp
/uSggcESBWI9z6stUg48FtFQHvT1vdk+5piQnbt/+7LGCnQGRvYaiRUxmie6MrFzrQp7WbRn/e71
DKFQw8pDm/5Zh6W0FtdV3RNDihCb1/UFPWySNzmKnUoun1ZMd7Jv571K6/XwoZWr1dBAICOnRrHp
5aBTgq/GhTNDUuUzaU1U7ok92LiTaXBDrx4/PTg+9eilLoCdcx7k64UgwNzhIM+goK5mYWzHCMCm
j7Grln8CssgzBtIiTkE5qeI3HZjJexttdQyYXWPHQC4ryqVfY+tDYqyaSScB1DJ7SJCz4UOHvd/p
FUxIf3N3O4F2ywbOEL5CwgQyQhJ/boUMV/m7jeZMo7u41ELVgyBe7wJG/ct145zOGbERuYeyZ34I
G3rMCphJTWVlItU13KIsFzVGo9greTTvQT04tvKTEra0dqmNhUi0vAqcbbGWUNrGQhP4GDYa6czK
M7/9ckMJP/o0VqPQ/Hw55RtNlSODaOKz9ZHsBb45NmJj2ZntdCEbfXPRxuNFPqdKoCyA82LWFlzX
xcd68xXnMB1xi9QQq3HETtcTqawW+p/C5z7PxSoVjM2dcosaGi5Cb+40yQSsyvnust74M+4eO4MS
S5tq0Fk2U1Ide3lKQWnZLHm3nf8bN6xzQmZT9hewqkNOOVFIZY+1E4h/K5EpKsULWecsLl28X64X
e6aAxjTxtqan6i3Xc6eKoHBwgxVkE/V7JyOieVSxLOASdsw5bCIICBA9hSFuK0bNh6g0729Ic398
NeFSADYit9B+vBjnxaIJZTrCgxs3QyFrqbthCvhpSOCAn2ze730EhefK0ZMGEdS2vxNTovORWB7t
luTSnkctDNo8tnPDjdbhFsgJWqGsnAlF1Ck+TRB87/n2K+RBeuho6VAsRJsDFfd3KOa0TzEOuFIR
a+tsh+WoFMDOMGW8CHx02Q9axO/jmrOe9WpFpYhBOI3cloW1e5J5b4LLmTPoeKm4C93VirNfce/7
1ZIYzDRBsc3YmWMrFbcKwVjw9Dw5Mr86NGfdKlOCuzOKGQlitbwuMIgfNsBeOxWb8pKw7Q5R7htD
+W5R7rWwGgn0hl7jtA4Er5muO0e0uiHA3zJC3xs87DzXz9VpA3viobv1qvQoZ9uOn+X9ShD0efnO
MvUGW/xGSeuMGPcKcynaJh6QDdi26p9svDnLXWbx/eXG0EKIpHhKmDlw0rxOur1S95HdUHodcfin
eRzhmcepKhv4VrM8oLenh/SuE94fbQWrtuHaOvBDDizVX+72W8+Xmx7JDCVNaeSG5lmoHZ73ISRf
3zcnrQhFr4YqVUa819mxDREq2SzmNRIT3CWnPY916U/yraQJVL4jskA70U0IH7eyy67tdjdbXvMx
41qIC+NieUW7NL+b8KaJ9dCc9D1x7AfTOlJoq8q/RbEtzlPfH4mUF8b/H7Nyie2aXzAA9PXmw+4e
HncE6DsREF4N8tZov6U2CJ9s14hlMdXnxG+o3Q2sKY6WltZ5QYavW+O9F+Jk/NyVCiVjFuXxb/1y
lIygOXoz5Z+TlJ5EvABb6XumJARQzAPzj5b47sV+gGZYI6ZhDKduq7VfkwxQLsOo3CaQaipcaC0W
FfIZSfEIwwkjTnHXT9fShRKS1yOlFOIm7G6rcr3ate1MtTdkAM6VhPoO1UioWZhaWLIzHB3Qc3Cy
G4f62F17iWg1n8ETAD+pz3VkCpqdd/LVx6jX8SPWLRqU7KU5UjNVgtrtKGIJhYKz4TSTN+lCcq2Y
oIt+RG16guDNo7F8V/DF1gArLczKCknBts8Y1tTSELP1wskSEsPKl2K5DPYOVW11ByQd5JNIi4HJ
2qoOwVJx3D69tOSR3GtIJfMCVniGFgUy9ZOBpgtN8FS9GFZFD5YT31/vWsC+883sCCqRQLXHRuK7
IP2KDV3MvYrfZfyLCo/z2lcNJReT3M4r0S8ba/xU0Lq7+xqspknXJOPHdsURHO13o6/buggVoxjQ
zaVZfVQhN+3L1OKpqNGgLa2QijkSTCgcTPBd8LXETi4Pp5taYoHIEDvu6CQJ/f8bDcMo0HiN3uz+
d5aX2p/+d/2Anbv+gaFFMj6ODCr5uxX4gOHjgUeY0Cb0bM8JzNgD4jCpRybREP6rlYViXq/23JqO
mR/eN0iqQI0D81JtT1503YUF6wIPM3kfYwgiIPQBcF2L4QU23eE8luo0ebMT9ge9SOq1FN10Q2iR
k22fkU4tDrRia0Ey/Js8ax8rXUdn7rB7oJum9FI5tQ3U7FKo/x4gL28WqhxlQDH0XH0hWRILqCwE
9snm6hS8xJD/2EdVTEsvshHsrFZt7HBcvNPlWXoXlTH0ceupNuDSPmON77c7k/W7CEPXWvtXuj7V
BleatT2c3hLxD8GsKiQ/HgNXOqpPzhWH8zapUV5JC+tES2x9jWiu9Zu8ngqWbrfeuttW7jFXYUaK
utkI02Kckw2ofBmppoICV4237/Qvom8MM+OKbNKm2kQTliJsM1zLQZHHSpr6BSpZWao+7cNwGFAm
0H6nkDmhxYsK1VX4oEpsxohbURD7ifi4gbs/RWpZDnBfAcS7ZPcF5wMZWR0ymTZSWynf/yd0Bz5g
QhoyMydK6q55UUCoVVgnmcByCEhqP1jxXBFb1ROywPMhWguBHXLcp7FDzm+gzfF8EwzFRyJ3IiP1
e8yXDCMkBBMz2hvBYYoaZeRRgSFxzBCPbclWKOJ/iaijbL1uASfjbhbsIki3a958JMQVxFUwnYxk
J4VJvEQfDcbiu/gWfPAO8r+W1renMBoZkMt1903Op4QMfEd73fFWXV/NjsbQ4T3eEUg1D4K99M7D
Rf4k6W/VdVlfNXThvDnrdsN2cZ3oh/BTyGMx9fGjwiGdIN5NK485KJTL2C5lG4AniQ6lpS0GkkEP
naSzShgIVjzJcTfbvS4J8x671YI50S8gAJlaFbn9EQdXGsOPXKZDOh8yEvYgYk2pZQP+oJD5tc9T
raC3u9n4hV1WHqFtBGbcDX80pmeiDswkYC6pS6djxwem2s3igt4BhMGa+DKvsALNiPOMMibxA+ni
Hg2aBF/HCSsceGpkciY8V4mlNNj+DKf38lCfzF+hMDOMxbC2mvAGxCMs6j++GEF/Es/s1TSV/1zz
DYKF8v0glU+IYE8tlYGpuI7w9p1sAl2ciLhMSAvrmUXmzVMSRNSelzV8dIO9JsIH/KbcxkMVD3oO
5xN4vFeQAcAQ76W/LT2uYs/7MBybEwXKl4ZD3CG8iWnPAIjJdJpGQK/nxwyt+kcqcZuwPoK6SYmf
JbMny4cwpHVXsqYa5/H2rSAF+8Ccl+FP7h9HOePzSwqt+NiP3rXeSGqsg8Wf4gAMSOn8f4hoTDcw
/7nQ4WQujLsG+4sUDBhTEDbRGleMJpDcBawwLJVJNcIOR1+djvzyWYis3pB/pUeS10oTiIYJQ1Iw
ciTTK9ZZU2vQaE4uipsf6Tw7IClpK1e4ya+o9Fnq3mDQEJKlJBWZURJHywqt5d7KsVyArdCAN1SY
HWFYxRGIS+S0h1TWNZpGnpVmg8tCQ4/3lSIW6QacCpz/2Uu+nWMD+UfNoaXqyTfVj/ChRQQCE4gm
SH0T+fpKjo4bmiHub/4zF6ajHuDLU1Wnk7gNhdgjmqDLQRyg1Cs2QL0NgYxlRzoyUCLgG1uJsT9f
9bteqjMY1g9b0YTiqHt3pp9frzWbhffazQMwVx+/ZIPuPMHFbae/hiuINEFwKH3KlVuDemiw8pjv
i774U5JOoduAE2MKkTAfabVZ4CXLvfA9dPUKbCvYKlxxuPLNSizovB/q6Nf0lyI6DMto9wsqvbG8
iT7KOrK8lgy1gwjW9DON0wCpBiCcM2IwLu7B7G6iPDCSik/blURjzYuPYB5/xSckcQGw/2wE1ZYm
kbFyBLcg7IJh3B8b2Q+wsKjYBbJKGpiSn/mRPnX34DlKsu9bj51Cu8z7t3pmM82ARjS5TjgxgSU/
y39GZT2tL0oYS8xmHgPS+Y7eAUbXWAFXrZONnSxaox40rB3/rBuz70rS54//On0MQKEdxASDnqn7
ne37DeNXVm/a5W8/fjY85HOt496UhY+Z5rKYkMLqsQoP7j4fiiXTlCAJSmOAEfVszU5eYIK+SyQc
VkDtAvV7OddaX311/G3fnARkzwLrSgWVHNxGJJjRN8W+uO83gsESYzRWjTovWYI+N6OVXcCVbA5o
+Hk9/MTbfVHCQQQH2qy5cDzUE+CdZ/rBFhfUhl30yy3el8NHaa1jUSpQXRw9AVqbKh5HPm6SnKOn
o3HqkBv6DBL1Lw+0drtEiFGPvseWXhNMJY426G24TRf9OyY1qPVL1+whM6OZbYhSz9rRD+icFRsq
MR9DHHSsiiutSMxggWcuAB+sNy2Tdue18JW1uGoEEfDxdxHQA/zqaPjgmFS2Ur215JPNuduhXeXD
PCHT0BUzmbB+ekEQBlHZb4Uj0ejYKbU2h/xIzfaW6ILvJr7/KwjKsFnGNBZ9ZlnCXBnzyVriHLU0
FoJIakpNbrXo4yNosx9VTqKe+/0l74kaL8vt1CEmLNlV0J4C1O/zIw5MAEjRu+372BZ/QLrCeOdo
0aWkU0293boUPeasDuUjT9Wx9NdgH4zYSa3PKmArRVe0nUVaRib5UZu3mYYQYx+D15v3dFxXKeI3
5IbTbPP8AD2KVBL5hwAabd3Ak2MgHLfrWI5nve/dRTDs3eXvLKC0Stg9LFqvBD53hMoqhiP5CHfK
TFrRnASWvdu9xfG72Qa1BOUpdR/MXZYnyNGzU/I8W6NOI8kk4PqNtQIH9ZDRrnK+cSrXXBV7qCrQ
254bWFcW5WpMd3IhHQ/dAAcOpS2V3w6JgVAA8NbdrSCvyLXwEmR6sbUqLBmftPpniIxoa/jP81VU
vpvmHU3gr9rd8R2YW4Otredl0NBXsT8kPa9yNa7RG9KDIDBNvRdh65OKy/M1X5INhmD9WGlvY9/j
e0gakaJqZOzm6ih5evGjM1dzZKwRABXB7FO77YshDIL4SK2tREqBjyZdhGOHEO6BcCNKhBj5tN39
k7hnlUp6MWghKq+ggff1gk3Qw17G0J9slFRoKMQs/VNGk1CfhKKnAG9EO7iszcBhKArJdkIjUH07
DmNNLRAnBDtIjrlH7vHeQymcwjpcqVUNvavvSjJPQVES7hI3UWEjhUBcX+ZfCfidNyT06COZ7QuA
zDAxd8ToNyrZ0cxIjxYtgL6jM12bw/UrzwGa2M7ClxfGSz+pNj0w9Q2BFTbzEv1BplRkoX8e5e63
0ixUJ4FQNkPRg3po5z4ovGbnFNxK2Q7xX1T1PT2cDnM81OSsQHOFbx1TO6QAKb372yo3JIpgeefw
1+0fYoD6kpj+RsLgAXfqap526XYQSFMa3aCIPJL/TSQL3n3yEH15fiAk5iSWo0HbTF1igPWnd7Yz
iw9dnCGF4vxa0rvGfKza82sDp1FHjhMhOrMjGEFb3kaQfC8+MiUbD+YEWIf1a4m3mZUsUSh5Eo97
off+XiXOM7Kiduc2Wn8mRudy29j1IJmCbaOvLOamqGijirzWVFcE5zPp5R2OI3K0GJ5Smr4PCmra
SuIp8VJd5wU8s5+YkcQUb8MkBkY+3W2n12GOjdQds7dz90MZmprkmxtm3vzxWcjE625hg1NCm89e
Q8FrhHAkFdVb9ZQY8rbVJQypUBosID/IrUNrv4LrRPrJD+0/byG0wn4ALpxVUiyeko4woxxWJ/Mp
lHlJ6HcnR3GBq4W1hFcws88DLxCXozQ8ma/xHyir2Oo7z5wovMb3/Q9COtUeGuqCDIPYmRkhJK/5
bYQAmP1N6xcLg3PnW+aT5aIZYSUImnfVdEfrGaLM4KWicvrxdhgz4pBxXWQnj3MU8KAOiZyUWqpa
BPReh1NLkPs0BD8fKC0Vs1N52j3yAfHaGx8tk/eiqEF4b9aOovuWFNl6TTxS9XQmhkZGNIBG2luS
WjOw9UtlUJNNNegx1LhFPov4MtKM6qy1S1Tkce4YN8AlU0Bfg+FDyIWuWT3Za8gjWe9ogt9ReHpG
A/DpHd7kAeHYzazeBNPncWCtrlKQ4jIrTpb0FfRX4S4aby2YvhJzstF9HCanUqvFBOEY0CDoyevy
Wo7DgXz3VkJKJhmO3oInzM0H59rAqECvbFL2aujgLVesBZynwoTInDllBWzfi1oUUIz7L53YJ+jO
jgZwm0AEcAbnenrH388BSrDktQWQ7oLwoU3IRfG+oVj2/yA8gJEtUaHSRZWsJ8UtIn6+Fihjh6N4
qMwlxQg77oIKyzvbOF7EiVZn8iywuW+u9J6zVavFpVuztm5dAD0KbziP9co82xdFWyQnndPuyQ+K
jrUNU5H6JwG2WhSaCPQpT2x/+pfvHdJpYUNWqll+rAkdMzg+Rka3YSeZuL1SNheL6IYqrFWFfCR+
scEhfdrTlu/uUpwseaBTzKAQ/2Hq8iyJvDa9rjnD48qoOoZMjNjA26RJCwmLXGXVsxQCWZ8OnUNA
2baNS2lUB+0RpAG1tg317LaNXEQSyfXe5ZxXYT4x8Dm5Cnfa5mGAVE++dnHbT7ANclOEBl4kjkV+
HH9YeSU8e2E5CGcHaMgMNNFd2R9YSQI7n3mFU6ZbsMrEmLfMAU9tXDVNGnAtWaW7+TQd02gSj5/+
kUZG5RnfL/i+A2bHUk1rXJTkV5Aw6C9BWFi0AgT7zJnobbivhIBb/WFNNxbbsLJYzQuMO1gt8kfX
2JCCMuBaWd5t0unI3/j9uKHJUBuH1EVDFWei8Lrd7iFmO3Hvey0UM3fbw2VxuTNVVtr23/SL/ZLO
sVDCKDFGF49gsyOgMtxOdHhLv5UBmPoIZjCX3VB7giZ8+H0iNQecFazrnh5u7mDLwsynsav9Kh/2
lOnp0ekI7hwakyl3Ycbrr8BcCn0YLjn6a/RtsbNL5iZOwqbdbF9/h41KHQmHVVEkhpeaVHr/imUE
+dyIxtHmkVu7t+TPIp6+775KLCKwmG/ZAZVjVWPJSdznVfabXr/Sv/UqsmziftnyxA1JM9JoDeiI
TCCJaO9X+HG4QbuDNS5ftwnL4xxQtrd4x+HKT9D7ygHVESALgTUKtFQm4Dc8g4KPk0rTrPMLi0nG
n/5/yXBlT33mGUtpVMzSDw0z5NHOm7ClZsAZ/Ws5vGYzdFRto6MaUYzE09SeYMGdB2udehOMt6OL
0vHXoRjIYpTQxTjbvQDmNI//G6bYBqDFVeHaJzi1cTumGRDzr1zPc5JbJeXtT8tF8rF72PKp3Wmc
7oUIMYHCBhKMVz/erOGWtvFJ2wUFo7QZQ2EWsTT2bGC18JJNOXS+8gq32QN0/DSMqMCUsPfx5I8O
wcrEWSVjBH9t3npt0my+lcpJH2FFq961heqz8QFhMM/mQxjWhn6pGU40EwBEGIFH1E0Ew7Lhv/J/
yf7TMrXJ+XvmHmU2MTBvgQVGUp+J1bibKvjYm/HPhGr5q3Rv/APK/FVL/rREqCn3qYuzSq/yM3of
ZOXQIiTzU/ZMnPGMXbvYAL8NUNTmTdUrIulzGv6MJde75tkOc0zWBODfx2vnhX8hUhfuG+U6lUfC
EfzBuqhpBLSShvR5I8EW28jwZz7tD8itF9eeaJJd6L7oxluPexppshFsPmKFDOV2vDmqtUh2kX49
QgsHZNTGRqTx6IcS6hnPTgZ8n2m77IgAisGAgtQjOiqD43dK1ZQh08l+cinsGB39LOgeXMUgBSO7
vDcJgu9bcMlcYopoJjBRC7uvrzva9JF/ZK6vGJZ4LiMlO6dOSD4qQHKoKQ652mwo/qJXgBGCPagt
cyxgeYNkuvuv8df/AnXHZZawfEatmLVpiN7l3fMhK74wSaxbJlGkhg/GvXObtwiPX4yVzvDe+71T
j4aSqKIMg6l9MCH1IR/mxTUEz09NQR50HbaDqHWAciPABUYjpBWr3jmY5GzDWdi7xOmxSJxvBTYb
5mdsAtEaJcyHOAlnKLDBkTNeJ75sjA+E9BdWqYKsHxPDgeBJ+KsV+BBxD07dxU31k1J9u1MMK9DN
EEUEfkYCeApe7Qqf8xWHIJHl3rZatJ3RkJ50w2eRoDXcXtkWqYqmiACFSpdatmtcm1FEfTlMCxnd
jXYRE8TxfJS7AYhcaB+WLK/8874BH70H8oQt/VHmW6rwo3pqF80fygQcnA4GVm0G/KgD1xPTmiT9
7o7AwvR1vy02TAAvuj2UfskBV3vTzONK+IFErLZ/WhlIwLrOvdlGJlrlIHtLj1nQehB5RoUPdFZQ
Niq+Zvb1s9qrQnazvbrxsaqoKRYwRdZxgBebsNqVbWGOfJORoCgiIeIQqzpDW+dK6YGZHO+XHOno
St6hj42uQOc70ygFdqVDx7Mizw2z69izYDK+7A7DiDcm4MCoYWlBhDmuTDoo4pAPS8y5+WeQVosr
zPy+vq4/0tDyIAxrAPhOb8MEsA5Y4SfeELLKz+2FJI773XkgQ5c8KkyscGffqEUx5Yc3TrZ9eYCF
G2bZm01ncVkcf6iKoNxBnYJyZ+HI/XkbmZ10osm2JXmN5wlZ7NsAysRhZhdB3qa0748jVjbWbpTO
vb9j7jWkki/yUH0Ck2pQD3upuuXexOxNDvvXyrv0LHz8rEBW9GnOy+v6iNJ/EaDQnH4Df72/wYvL
nh4oDWbECgE1Mb3cNtECUUzVZbfStZBZB5txZp9orI7D34gYUBUseodm26W9Zf0rXGjV6isyefam
VLQ3cueb131IwcluP5jhwUR//4UDxthsTuqazAXH6nXbArOM2cwcBm6E7Er5IB9O0xweHkl40YNc
G3rsGWqBfs1hO2gujSxDU7up2quGVnW8kFDkE8cNbnVrvCE1uSDTFw04wcNFKZWuwBF8dfRJ2ktM
ghRBzhsaZ4frb10Fnb5LSZk9rD0D85agtADbBorI6uQgkpu8I0bPNz8+8DfkwkH0gOiMIcB8m3Lt
1ppuZhOTuCAT49f3a8W+ORoryVfEBCUGpsuxNEzf5Mz55s08ByymXUfpY9RxWnDvt4VNcPn5u0c1
iVEmRjSXLHKf8lNKneE5/Chi6N9t3aPxba8vk1ly3W54lScj8b0lDKnYCTSZ1Ktz7CZPogeU496K
PfDyO8gKtkF3EOZ77OM76mEtaXYQANoIhhCnthLfcJWSlVkOptIplALjnxXsLVKhE4ur+IYgvQQr
5tbag3C5SFRYNfJHBdWjkyIMsQti+oYQmljUXnpO00g9mGsTKCCzK9CfVwnUAlRF8LQKFmhB5vNx
9aLDp6C+AZ/DZsUGuGkxpzE36VQ4OVOeG5a91Q/0GwYYtKRoVD1/bNH4YYJm+2M04mwV3G1My+4n
P2+w21gNG91q/4V7DHL2FAvLZRYMp0MLJuVYEJy/Uc7dsXzJe6owIF5tQ28FbY5J7bCzcpkCL3eT
9I6w1fDHr3PfuetbGPmhOdYrGvqHUSKvMg1AQxMd5SmW8GavKqpaw2su0jMYV7b8u1Q+JUT33eww
8SWVY2WzFLB0r0Ifev4OeznrXg9tgkmGTf6JerulX5wgugKykfLb/RI6TP5eCzEk7PAORNWxEf5T
AUht733ImLcyf5NvotLPx4DbsIoi40C+nh6cfvqA8onk0IBlZR12GVpZ1S5i+O66wuD51EY7ymbR
PoW88Avi3b6tR/8Q0UkirhDAM1OeOIulfYFgrHKQpqrsWD1mRCJVYF4N3mHjc/DiyapaBIm59IbJ
mRgiNAdI9iAkZApvIffH9iBQJj6H1HaXj2vQkJMjmYm8QYak5NJkOcSIBhJ6RhHVI3qb2B8PIQCC
UNDQWzlgxkqW+xeNQTer6dIMFCfc+dRoX7AWeLy3ZeyPa3OU6Vy0ZX1twuW7upJkfrC0TlwOJdyT
/Fzp4hIjGSSad3QsI2Xlg1Ma3Qd5jUBU0cbTdwQiGPMSDDwXenksoPETo5XRistiTJOjyKQM5Ony
BQbyzPKEhbJW3yKIW3FocPIGgG5+z63eAf0WK4rp/UwrXjwZrecfgmca1ErrQWZzC6+MI/oC0Czz
9C8C0d4IADYJY6EFhKHRJzukZHX0y3isIJuIbMqqPVs8cZgSMgfS5o0a0NS9NLtPXcSCVH6XZBby
dlGjxluyOwx0Ub3woH/iWn7DueOj/z+5cx944xcKegiJAYZbf+sGmaMQLFUCCd3Le5fBCKPSB1nL
wlhxVda4Ga8nc7b8N3VJgnJCCFH2F3sp57lFdDl59UXN4zwB9AhEUZQf4nMoifl9KrufH9RqHW+2
XruCsHWjBmGAovkYvzZ3xwZAe1KdPjqNpvhjt0pyA0UY8/2ijNjJmB/Jhp3bWKjETr1gN+Aur4qS
zmX5XnyOCHA9xrpzlPaNw3y8T1/k1jSyv6/bD8Q7SBpjZag2F8zsScGdy1AmdvDmoyIHMPgj4m+L
U8M/sZHvaLI5Btu8ldsrMqd1049n77Wummx8GT2iQEWxJubCdwG2fqrwUAr/wi1xcT2WXbN9JMCf
v/ZF+7tFS1jdrgAhjhhWUbqw2IEdFhmQEkvUhYsHmkpn+My5NLO8TciaEGxYvSO6xmsODGnT3Dqx
0c+lDB7mc7tOH7Fo5XbgIoQuLHVh0nMWxKClQSBMcwXhrFJ+Rz1hx3Yr26bLjyrMQ3UqP0fkNMHz
fJ3lARP4aZGzAO+BpH7cNrpnQElFoZ8zo9cunLAd645bhpwbfDGk4/0BAPh6F6wegodHuh41YKAE
qxlZHr+8bBMM7QVCN5tRc5C9ohx8XzekpiTlgfgbnt0htfhQEjXY05XOGSCU+FFJ29w4Ahm82aSl
nlbjCcoMbjMDPJ80UfOGot0T6E0Vqh0jEt13WdBvlzcclZDTeJeTZ6UU+qVWqEpUUDY4juXzl5qp
WObjzIvHaS++wSoagUEcqE2jjOAGARExwlygvYWOGgseC4xZw8oRydc5Qgw/CP1jL6kdUiQlPO7G
YJ8GYIcpTDIoVpPXYVgvOqBocddlJpWjLUOxvln87GrjdTziDuhKZ2Vi1vgnjEEBuASjQtjKPNwQ
11PoZ+gtv2zgod/XTw7Gg4FZA8Tox9T9VQ23Nbi4Q00q3UrzvcGmIKuf/4ru4yC25hSrnf9PBE9O
5xPserJ9m6FbJgOV7CXXfqSpGKNxMlA/fTCaNCtiZ5CkDxLrry0ZRnN1AQ637p6Yqb0tt3cmzZbT
tjD15pIjL90vQJDIyefXEWNvYzK2f6fcDFkW+oJiV5hz+3/t1IOGlwQ3Zqyo0x9nCvD9wvM+s/mu
QHhyhFeRqKslbbRM5vHozpyBMY04ZwvcenyH4KRJV7eE6ryoOlqCw5FaXD/PXi1s1x8Y/rRr8JyZ
tDDkCBPvft6o6XUtBNjNv9oHTrj7NfIb+WMoPLxV70laEaZkFke8Hn5CitdUTch432pj2Qhff2rQ
DXVjXVzFX5K8IGwCuHxTxQOItxs86WlE7Rts4FqgaVCPXi9wtRtIWTIbjmad7SGgMzUNiC2ugaG+
CJEQumdmeGGoj0Kvx5RGcjvXYa9eSHPCf0UG1ynxyqZvC1ppqihFLnLBi0gYvBXwhJ3x9lpaKw8G
cIaGR+ZCtgDNZljZ4KyCg3/50Fpdl1FofqAhLRbPLRXTF2hPYJSjwuYzWxszuHoxRcA6gYOLhqvV
eZWivpzjNYCsW9ZDZiY1MgKrMmo1mkTovaiM1WuwAq/Owqp4CUzFV80V4d8T3ZfZw5h+PzixbZ5P
aZwwxAOXoLzY5LJsvyB8pMjIXoo34jephcCgLM9228rZdM487s3lpZoLkWXRxZ8KrOyVF7ESpBgT
rCGJoGGWQaT7b/UCjzcan+j0HGkhcUpJGNoS/EVWotsU29YdmR1eZ/PLn3pvKqkEVmqBilGJ0tOP
mRrNV9GYcnp5OPEkF6VIePDppni7i5IQJDU6Zd62Fmsx7SDP8GfUPqHf+2xCZ52DIPIFB4NKXNEG
+X9tGQh83PLS4zcYvjC3lxQhH6iYEQRyvHzgurGg0b2B8nyXlRaB/bch8MCZJnAEGBLvYjJ6u5Ft
ra0xU4K8sq7KtNUFeCP5NQE4POnGTiiLhA5kUIqYQ8L7u6TPfbU+MvobpTqGlvI2VCMtIVCVc5Tn
khPzUXj0s4TWJUxsLXStGgLG5b512M7iiRdldaB5PnJe8eeK5g1n32jFpaQ4NZDMCBPqlxnd6S2g
pe3wxnKmNISJh+WIHyclo2gkCXbni0J2x/TEU6gqYjuZyxpAj9fNsOpG8YIkzAkix0oejZ5EwYVf
fDfRW4PLyo/JzE2qPJYbFvdusNZ8uSlkIekUJQu2GkpC89loskzfufOrO9q42SCFO82YlB5d0NcS
gxIt+OTNpaNqkPiHJE0ZA4TtkkzF1rnmeIRW9W+HVZ2Ci3xsyAzIxWKl3Crp7ZB5XP+kZAiohfNW
nl7yzyUCI93+Kecw9EzMYbTveTBV6pcx8Oi5lLQEzb0wUJGBOBaSBxvBjmXeVHv1VBz2MNJlRzum
XVHVoSlkG5fSU8jmFw1oQborvfyetAMbKVxX1beNpMJ+Gg6mBhNjTaK6THgEvKLvdseukRIkoQl1
K80YNJrNPvcFrkmm3PLmTw/JjIIX9bTQfdbMVy5DnuYJ3JOfAZ3qQKrBHScsD/E2T1teZSDsySi7
3a1lFO2IyoVsN1wB0n1pyQGEEfCvRCyeXAJEHi9ZGHwdbIYCz1POSLdy1EvwyBP9aowO3AbyD6sv
S+kT58GuiZPWwZIS6ZKVG9VL/d6o4HtDkTcvUK50rPWqDdF7AwmWNnSK5MTGdED7ZZtiFoL+q6Nf
ZJuVzIW7+wNViLHA2yTskqMESBpRVKixnGtf15O+dhzg3GE6WjrjtM0/9QKa2YCsWQxlVyuSjb93
8UhDvsPzdyemniKuXHfsmAWeWjvuKp76oN90dyWN1pumOd10exnYW2Kq8zu2hYq1SJzccAh9Itvz
ZcOJRpk4zyuGDofF6XuAQk52aCnfL7urpZknRsV2+tcqd7QnLchDEs9onohETtc7N/tqN/Ppuwj6
KEcw0FbQOqEvcKVSKzcI8gQR/gxRzbRzxwnan1vhTBl6qjnEvLxnwqd8o+1lSlUj9BRSwtPJ6eVg
HS5PCpENO6v9+jL8GRPvRzbDxhiij0CYoGtsA/OXv+mzjug3nQ5khkC75jjQkfgtcm13N6PQc5sB
xd+K/xSMcYzfbT0RuiHojYjW3zIO4DIpOlmv5G8Xh7HYgoAbG9aAYUo2gEiP/rACrMWk2QXGaF8g
gsx+R8UuDQjcoA9uympmaTd8KzuYmDz3W12Wi/jIRqseSihhHQ7jMSuAWK3txCPNriPxy3y3I8V1
y8WXCPymOsVWItvN8CtCruQCeB4njbmEvPUdMlaqt2OrvtVg1DnbPNsnEL03CHNZjmjfqTx4ApeO
hoB773QMKHAEjv08jDHPkdLNvFp+wNIh/sX1n3QBMHxlb7C/DTTIA0lA+WA7pUXhU6rTB/7/MS1f
7ranEe9e4TVTH8NmVJa1kKtFbVgpYWSCb4r6XUkswbB6I/s9kC1zEDaOfxgrt03eZE8KAI2ul8wE
OME3I+0BuGxMIcL3XsVSWmUl7oGyeLl12fATIdEZOhTG26aTRS1heg5OeReqvTTwIhW05702dnhi
acB2xfXU1Dru7SUBWwZY/zQ0wp5rfrvzniVYwzHHJASyUBysbaJ+LNDqOIVZKx8kpsfnIp7MG9l2
uOP64jTn9vhf9qV1NFU01/bIzKszyVQyVVeAwdW0m4NGrhl/msAHW72qKfpY9CNx6Tp8wB8UnCjd
VVs/rIEsBXxDkvN0Q/vLcH5u+eBIn1mljKFQtt1K2FKt5GP2BNq6qHIJSMUooFA6dudHssbj3p0W
HFhqD7tZRs9HDanN97spU6tZJJvB7u1sWXTXurWXBcEuQdHDD5XUg6/bNa8WErABFEqv2VLE2ozm
0cI3J3A2z4xCQr09zwfNLjo/AfjJFei/EOD8bufwburIyLPiI/eFa759Pa9iC1PeX2vr2mBgWIm+
WX8LNmTdrjv6DoIEoxn4KcT3sYxC7+aT3JYwfa0JNuMcN3cowWVJx22759VYEaJtG+RXqKVrUnLZ
BzQAPMBqy0o7sG4FTns8cUnFXBKIvSv6AAetbgQL9k4xJqv9HjTiAczVNIJSp5BkCfSVTFhg0DNi
Q7YpHF/7YXIsPqn4z3QTbPJVan3UtjZbFrzhLJ1hqoYW6NdEMLcrhSmo4OzFtYLM7zFoPvWm0HCK
8D24SWHYpZCFp9i0w+GJJgBxa9ACEo3r/4KoYzPJL1qQopuFhJtyy0jflm4AibTGLrfapiiuLE7b
HI18FFd8q3Emzu19AW6v1apnyBIoMfEtt2Ky9wPwVH1Qah65ngEoQz18S8uVPsJPVzyc6CanLLuU
2xP0hkSbSAtxj7xUtgDHlckI1tPdEkMiX8JkUiaBH53AnlMW1dnzGNR3jpsVGCqC2kZUEbXRvUxA
rHxJ8GTqV+RddSX3p14AJljDT+m64TiJAv5f7/cWxiU5Tfpa7LF2ancydKD7QTGHOPjnM6dLpDkD
TsBPbRFDqeu7zjPohmHUYmeWJRW0JccQSLDWDV1J/TM2cMvRiWBhdFtNhH8hYA9uPSCC3q402sbh
5pNA5cFYFYBJqf3347gW4xJhHyWeNqDPmhS4Pn5sSkbh1bFr2zjdVFdtvdRBFo2npEUTogKLiWnB
UkomOezJ0StMKJgC4F6a1ozqlJhLCkNbdkNzaWflNkeX265dDAG5aBNm7fg32vyhAtLAe+7tdaLT
qR2bhE6zHOqbDm/3sx7BUfE+NdcueI7qd0Jhdbnmh/Hn4dSxonHUhTtptEG5i549WHQP1UDyZK88
nSh1IWpNxP3wMiXOGXrEQi5xnde02iLtG9aZFjDVh96Qi7VdYchyil+po2u99UpyEfqqZm6KSlQZ
j12FZTqaEJvlqF8dmNFng4zJSXXTMkjtSnXhXcU210HKRidmvdtv+vteFEGHfDdwtreDX3pDAe7o
VUmoA0/OjRJg70ArhJNEvrQSTU7U7/MAXLfHIsRTfPIl3ndh9DJgGbTwrY23BxB2se+2Ip7aHPY0
I1dMzsLqEWGGRiXF/WLgZQxrO89DOCJ0q8Xoi2OGC5HabyK7jAuMR9Rm9cpfR65HfzKDtAxwUwOi
1A4oDMz/riCB+fBfbGAXNY/Xye7lK3zWBqBCk8ubDce2J7e540IqmoQzunlZ6R3VmGJ0gDWsKigi
kEXU0+V4GzeIuSiO3OsFvSA/BzDEh2gM1YKpFUC9H/YuLJY5RIOm7GNg1u2IrmiQK0Fce20RrUxR
n6UXMzITbfu82Y7knmpyYOY1lddfUErlZpGNual/iZensmJCCkMpzj5uf9j01bLiS0c/4XbuX1Cr
zkKxigzkGwor2QbvhJlli0DRNg7McNWuSDgFvPDv5X5ADsNF4Q5Zyi1BWqDCaU+v/aeY1RsDabTx
rBUQ3SHEXPJJ3sXDcw1AVn5dhwMc6XnkiB8va0YSCFRDJvgiznGAmzAKyiSl4uk4SxXzGCVPeX06
rw7UkC0a2FJoKgtq/Zszd2OMEzvYMzq8p1ZA1x576l6S3bYZ3DFUEUvpykUDh8qVfDyJ0kdbXPt/
9M8uC/KnyLwox/l+HGCvkY76xgmzERtIn4z9JvHuLK4C6HTXaru6OvzuTix3qBvfzukQw6MKQ0LG
fGnIa8Si3rCTEZ3l2mAxSDwP/59hu7QgbjNwxCUqUW8LEEmwSXotg8LQt/agiD9DwBNzx7E9UGzx
kae1b+5sPF2SO3akR+cBZ35+MDR5kaKY4wphhihq6++pdbY/WCdVlHMnDiy790qNX5RiaF3Yejh4
QiuDwkS0YzC/4Gy9pTucpz9Gp6Rdpjv/0ZTmyZCHy9uAFqlk2iujRb8FW2g+Ewa4EC86Zhp0QSdx
mUvBlKQKpOguBLqKbEgxh+3GMWMQA26WKOe7YmRWVBeUn0BAudsKCdiMrV4ZC5wfhlOZbXnt3wsF
HTJ/f2HOj/ZFaTcHuCTcfDHH+33taA3DWQ4nu8FiDJCCWsC0+rum4Gd03R5+9NpTbGp7nP1vCC7Y
m9kNgcso9OeFhlkMsNtIKb6q774xEmPg839WgquOmtluNF7ViWq3Uw32uZWvQ81sOrCQl5UM/QWC
ggI2h+m+QBF7a0qOymVbLEkpLcLOuSSZVifEnulBw8Vb93S6+rCFO577tsrpDGK9DWejE+l+0s9+
1dL0Rd/+gpNZyrfido9WYnylhdiTeMtwVD7N9JlH5AW8Qjz1d83i3gdzSUfAzfVb/jzXptYPaq9S
iRr6QuYb4fdCa/xWfRZMvMb7Ia7A+8SWIO9Y5ezm6bd9PA5e/3T7AmZWV2BtAEjsaNbtu4DaT4Bw
paaHGwD42dqDFnbsGKjMfBtGnhodCm22HPYC4JV0c5Zx/NBLFJRkJeR0XA8vjwevgX0Un+pU8w/a
kJJL9HYF+dApPBCMpo+Rwdz0vO0QfA8qYUlLR9fo8qUVw0Jnj4L7Qg7VWWRCp2SfU+uuJLaf31qW
d8IOgnio499iRe+PgFHPEa7BPAuxtDSnVn5jPHm/r73EP/iuEoA9dP9RqpqBLzaKkw+qIfb2OUlN
I09PykxbTda9supR97Q42AoepBfsw6lOQbH64VCR2+EezoMeTvh70ccSvvHGJRRqo9qImhz0hd5M
O/NrYg42p3opl6vcaG+P5DrhXeRch+CvhkHQ/ShqTa6Uve+fFL+r7+SfWLED6BVh0uKFFKAVxziT
UndHE8p+YnckTHWipLqPPveWt/TajB3yXoR6SEf7b6u9u19yXyGHdME3t2fPyqqDReCQ5/KBJRkN
eilWs7PYeC21bih0VSWkC/r+n2DrHZhNE5kYmH6dYBiqxBTc2aRY6s96ZT8xaK8sfP4cZ63130nP
B2ohr6YQi6hdoRL25QVxqfmHlAkFsMbclSxLVjCDnWo29yOruDR3WotG5OQY8md1598jA1xz/0mv
EANod3LZYhErllgPZoLccgoFzUdxEAlOqvzDYfQJ4vklHcXVGdLR2sCcm0q2jgc7ZhCNqueOeMXw
5cJA08v4xajEjCW3G4sioQKRbjJt5gg3nCYVvJxyH/ZZuGhLEO/0bztH6mlkUcBMihEHchYuDWLc
C9CwcJzJVY+607kdD2FJO266PA9lPUTCzAwNVdqU6UYsV4XRkmEJcsJ0E4af0NTSs+ifnuWyZRS3
kdeKTac8e3yKTVqLGF+Vz1Jw9avY2/BZTOitSkR6CTaLw0tXHLKs16rAatTj2Yxk5P9KgcjidYoZ
9NKZnB3czgSCwNCivaUjGmEbFCw8hZKwqIhmdrGPJ/9wTSa1fZpo44QB/EdV90R7XN9hZn5wh5Vu
3zcEFq4O5k0gCy+IMtU0YyZ11P/vm8lUAyYpv38M62Xe88PJ6Gogc087kj1IsWqTQlTf3UvZLI/j
/IMdU7LnPrhh6qgf4t7PQNcZdE6e/rgOpOOOnALPsMNL3neLbvHp02yMvWR6GJzVy1m982QqwuIX
bFsoBeyLLpz1VcG1uFXeUnf8mhRDfnSGG8P8CXvoAtiPWPx6+Ez8YofCXIcfGHm8ESt85A8fopbz
4HucdN1BjZuu/WCwb8O7eILVRdy4TqjncS6UDruuvD25NO2Y2uCz470i0NY1gnavnhgvtP5zrHT6
sKmkO8IdOLNuE+Kt+/SBWlWWmQmRnaHSZNQ4vbq5GMH7z+t9Q1su7e+4qYX87VjrvMAWHtOZ6NlY
F+q2lUgPF4JFvZjUhGrNponpibV31Pd4nUjNb4GDbFKcg0R0dUImIUtQLb3HPqdxe2ZFdxL2X0uW
i2vHVAm4S5P3VYJ9L/2T3r0cYvuxzMe5COVUqIQFVxGm8fB1lJ4AIPc15KRxVPOVAAQY7pNgZfj7
pRnS/H+JagVd5LTmJ4jSQhTZGk+PK7yLb4rViiNQV7hAyESqG0JLfJ24LFIzUM325AnoeTkw//Ul
dKYwfUU/YDUQyH9M+UK62AALnkqWj6DLgpb8JWKc1JitUlk1zdARWxAaSoC0BCzDHL07TmUZrCsu
5US3TfnLM9NdGq/Tm0LkAdHFo5GCttKjwrbNoHSpgjhK+SF7PO0LBbC07JM4LuHCEmjrnFhP2JNv
0UeY8VS2sjsQBQAchvXoAhbbAj20yxuolkJ3BlszWh4E6BFbvxuki2temFynuU1E/LXemwbXfO/W
IGJpnDSqOjLjfC9uot0G0d/2PaI5oddK2mKa749XhS6vgATR/uwBc3MHUmqZGOlYXzdi4TlzQXWI
1DMHcM/DkNvD8YmhwGVRgGiuA1AUzg7ZuPqpkzrrqRQWsqoQjUSmGr9jDllK0+/ukrAAyl9BlXtb
T9hbLJfwt5x2db1HDLjMa3YNCPMooAPl738MweBRrMKYSmqBqso/AKGjM3pfxyBjrP+qqPm7iLWc
I4rQ2k3cFRFETfsQdjbTgkKFVTPTymrhj6COYYHaBOc/H0VyXLFMY+Y52yoWwZ2sJEqo7Te4HcIZ
+1g9V2Wg8NycUXc2MJ+4XEND8B+U0fpp7u77CqoEoTcfNgRpEW86dOMb3E+PgTx2RpE3+Pr/Qxhp
l1jl5zdf7Xd9Ub7PraInQLhYQc7wN+Gx8NmTy0et1fL80UBJyz0OxKRiai3OTJByzV7rJ3PRTcyp
ooQGS+7IUdfRWKoo8H9/TE+kzbOwwjrfspqNrByoNh6i6NINlltknR9tKVZdP2Ie8Wmjpvbr1xdR
zje9x/cX3LkoHIPl4zSOni14cwdDUNtPnTWK0b2JMbpG0mqcuPH6mx4+s1PnGE1g3ulst+AL+WkE
0i/aP0so+GqCr/xQ5fBB5RdJjTiuKxTB2ZeOxHUG1cXN9GlVoH4cQW/M3u00l71BFNi/LY18oMFh
k3ibDtSgYvCsZk88mdCZTHwxsIMDooKUDekhHFQr91XDzfhtmcr8FTXVv65rLdrKfKV8UEesHPD3
t2mGbOadxzgpqpwSJsMZc1pl3o2knEeHPw7DTS2S43uWVQBwHYI7vMO6eeAHyRYDE3Q56YzwTrN/
8QvFTzWyZMlHn1g4iX3vTek9kWYOYsgyfSWnl0sXlibTeeXnuAvcAUFgwjiVjlbWbFKA8sDdEPls
YJc7z3zrCkugx3uyQCY1nuTXQKZg55f/MaY/ZBcISjVscytigB1hvmIgfG2viaRpXwuhV6whyt8y
jtyMyPFpaDu6cDTMFe45Qpqh/f0wh+Hg/MxOVfFFy0T14e3w33XaACqI2eec9nh9RN4SYhWOMO+A
WU6/90tz+zCo0oS0irJn5bLfF61bCTehaHkgb0kBHN5fw20o31KaIUFCvd+FvToa1tiUzpiNnc8W
1dLYRqdrTEfS4wc2IovuQFg3GaRUXyEJoaptEV04iMrYfOlqffhhTETEDzj5NVkGmRpU93gWLyMk
ndcp1cnt/c2T3rI6zWE5g0LQ0ST9FYpvwfrjWxAiVDrRyiLKb3eMDMFNbHGr7wtiMJ6Y/5RtC3ne
UCL/YZsdVZvBaW9SPw3aue6iiVK2+DUuQ2zUUEYI+BVeSyrOzohM/DERPy4MosXQ6/0AZItmEwUe
zevtfDAVsfFJ6W7P7slyzG0VSELuyxVr5ftp6SgV9aFdCdctX+Qs7j1SuiHfBYJt06DZotaOPMyU
3JjqOtKHWlN+TdoBLXjW56S0vzlY6fqvkV1fiz+Qnz89KQUbdHQJBM1E+1ei03itTpSsMl28vrWX
3MMhpIXO3+95Z5lByCA5zy8LQSQiLi4gmkvAhVLX8DvnP6vyK/IpZcKM099hzVWdwG7x8ZWEQn97
+4Rx/mZ88FQ/nYZtlbC5LqAQXSTCD5VHBP947LrgJK5QfvEtHiVC4XxsIzMP3vtZT6pLSMRvNGxz
ZMgCBeUdrD0XO6BYLJf1k0HyLwfJN0mPRZMdEz6x3z92SZf0PbgNvbtsyzKzqcdFLSUtlSJMVEe7
EIlGqeOqIKgGrnAEykpLcDDIcfsxQCq0nMJ1fz2HK/ysl+8Up5nOMNhzbuEqKLUWpN5qsjyBuiTa
YkENHfig+lw6CFKSeeTUvI8OaRx5jysVaMd4GlhTw7IQ+owJfI7lk+NfKMYVQ3okuAbboYwX2Bmv
TN+ED4jXtKqdBDX3l+S+U4Q48uliVKxq+HXU3evoxk5JWgip5kwJUs3vIWCLEf5mkhLCNEqEER5W
46ZpBsUPDLPR5/dBuNAQLm46otNENFPEzESDt1IKQ6uHwFnpiw+Tp0/bWRExMwS2c/vZdksrtEnT
ojlS9Uha5QQ6dRGgKSARsavcMCqrzWeMs/bPu9ATFduBUqOlXjuXIxT4Y6yMpCOxkuBR2+jATsko
2AdpvqkGzpzq/Qe5BUmcqACAf+VD0OiMwPkDXzSKt4UA5bSHyJpKpEstpmIGTJBATyYX1AZ0jXA1
OCkKVjoZ4ISr5JSVDEHAAzFYqrE8hyyGb1vBnIu4zkiEeIfC73bqtRfBmz2hbBI4Q0GYna9Q8BXw
9wQxX3nW3Zr42xWFIlDvk4S6yjp6qf6AXe83CqwtR5J6nQfbmm8xatKduYQVIRVxPfCN8rDDhnAe
kqvG4NpppA+1r6MI8xfYs2sFQwnjUgFM2YV7yy2ElYBhtiSKPYtf9kyMzx78SCGXHRgslGvgHNyr
UJttHyE8sbhyVUYYq15JKYGihxWlvwFece/eTjGP8Ejrz9wuP/TLVvA0J788kr+InqA5uUNVmnYZ
ZaEFKGhsIjAw6b7FhG+G6uPLsAusSdZtstHB/hzdLnbn3w4Aq5chZcXu5l5VPdz7KpYKTh5jzaAI
PpYlmzW5iiHoJdE1hyP6J/P4hW+tMKtiRCY83tSnvIUWn63KnIC8NHf1vOXzLfTJtshYE4uylUAz
OiI85Anxf2QCC+D0TzLcEtgy7sRQbPTMORZG9EDYIAp8Bj/yFFqYSKWT1XFjZz52ho1NB+YD1SD0
TMAqT7hbyKef3Snkj0QrlGMfoLklmCyGJFZt58WhuuTMwCVVSzZVC1v4cIPvJtZF/dYKBwkXrYRL
630ocnkXAvL3pJQuIBs1RH/VdPuIc8E9rzx3YjjZT/jyceN+raxCbb4PC+j6fFDcDn5U23dQ6bBJ
1ug4iwTZblljATUmf8okwhSXPCqlU+sGbHd9tkzALLgHVZjyaxkZ29ULhnvRoZmEuPgFhbCfIYIS
MwyjUVnnTZHbsvyGt0ssQDVkcEV18jJJnbjtSAwd02s6csoHLC0l03HkNEiMI6BKq6PrA6NVJGv8
VDrbhs3JFJw7FxE69KZFGXZpA6O7B9A3NAGSS6ItfTd5zdQW168DaBvGhB4aYa9kurQDWZNNCaKJ
uFsnz23ewPXSIo27XRA95b9od3pawMiSI5/nTwybB8Ca76iQDQgo3QCwjRduZGnthkW/xJ/idHzM
MULWjWChlRdRIqfxlf373QILxLfoOz7d9nJ3FPCx1S617nJLkWaA1YdnHFFCfGt9f2GafcWXl8Iu
GEP8JBuRSJJpIlvjVrSdC5Htfqc9HYKAxWBlt/YECDkxu6GkXMIzZSsTMbwhKeAe8kLuBw2lmOFS
XpNXNB2P8q2wWy5NPaPwjvOxAaVW3Dmnexu3LtNW7oD7NN9HTgTb5CQXfIoMaV6sy5gc/3i05jMc
UoBfiRJKOEXWgTcGgDTiFLNCpZZfHS4wjIwhZD4OLMmVPd1JsdGlD3BHHuVgtkhJSwg4jURrSLTy
1qet5yJov+Sg7By4EIS9Ag8LOElRT9gvumUpvwwagWEYg1nYI0ZNJN+ujLFKPiC+PWwvqAgymV5u
mwoHscBxNumOVNo1wIihOFVnyZU6TGSnRQNv1dLDT7SUQsLV0UoXgSx0e1sltKqMkdhCKo0REss2
KivXBBeJte/bZ49KDHuQB77X3Q8IXj908dcsTdkXoLI6cKQWcyZ68o9tOe0JKfcJMtUjZOcjUTkZ
5vWvdAeUKnghAT8pnK7X5KUKuBjVFfSu/mKVepyrPVtk01z4Onhz5ErQGRBXZFC5t5xA3ZnE92o7
6KQfeJqxGH81kRe0cCffJIy4GQEfNHPy6MLCue24lEyv7P4ZofCY0z09C3FX8pkZUtEDJBYD9Taw
w2h7ZcJsgSt2mnIyRsIgtev49O05S//srcDB3O2wSPjLYy2Gqlomep2k5BcXavWcZZ/mEyKm29NW
2g5MhXsf7sVt2dHJA3KSiGZBZ+zcobFPsmWHhikagPEsIAnEW+EfG/XvPLuzMDpgKzkdbfCysbQU
2F612E2k4/je0LsklfhG9DruGBlZok/P2/lq3GOo2AWPg3qtf/EoPKNqnIa4aYpiP5bdP7X4DZIR
liK1jq1bvqX/r7ujrN9htypw8gNBNg5OHeLRG4ntt2+JqkK0zE1upPbXDDY8Kz7eySWKn4vqyOtc
VXjvVoPSEjPXx5wDyDi9nAYQvO+PTRetl8cV+ccKxPZ5c6uqC0ea0HcyV8RoFztivwgO9i4UWbrv
YeG95t+3Cv12IedeTw2k124n4lt/zUodhLMEz1AAB/kEJMSru7rvT51uM/8myjz4OW1cAA4t9562
S4tDZqiJOF5VFE3EHT24J4/4TxrFe7y0TyYxWbY23OCb75wpOQ6HMj8crV5DPMEKTGF79RxGJ7kv
X39ZeG7khB1oVULFKhjejTLfHg+6nE0MJv/IL+IAk10JacU1VkyyhcTL4dCLS5TizXTwfmjFQ47R
+u4Ih4boe60kCdfJCT5pA1BYaz4/V4V0BVfxtArSSivPYn/yNO3bX+WryCIVKirY7QbNFDA2s17A
T6MYGgFJ39i7L/CE9rEipgzvB8afG8FoSOMg+YBASWcXrzXiDpkRI+GgYn4YiP4qysfUAroWNQMH
fAEZEIOhR2/FtxtpCeNjvXywSKNDcCKp/BvKIQwRiXZQMUSgegi929IyQBs9Av93W6owGeVLHLyh
BVtcpCLYmKHpjuTrn1Z5pCer9pcnT6TDVg42YC9gAwiBB4Z4P4i63ZR6fCNxvc459RAAQs+biaYc
MSCt1OZmMgPf3xrAJkx6Jdyez5gTjPXwCln2tTc3hZ2Rgi+fYWdH84HkcNa1rQgnBrV5A7RDige7
680XY1pM4IHHJwSm/nC/62YWJLhJzCz0HLGLm9gm/EDGpXwyfJH0CaJDVsuXr3D1kt00ATjFLUPH
ofYvvat6qsZfmJymqhtYn1uslFi7t/+kyjTicCrq2jsWURNtEkqkM2tPujF1T7BtFgqxHbae1Hbe
ugJ5/xp+BbgiGDpT9TfnQ2AMZ2lOZ0bdo4W5LRmP2Nl9lxJigQYTfqtVCoj7+aSJNEgFggf3xj1K
b5E11ueEu9qYmJrZWArR96OLau2tlqAfRkJCtlG0IGdLDNJKas1/lDLGqElfw3HzFtNCE5ZCs/B7
5YGDmkFLtuvumykQCGIiDHxrxp8kn94LVRSXNG75zctBhtUv65YdBv0taetPW9v5H5D/TJm/3APf
QnADH9LJCoSr2Hetb2BQirMw4s1nxJLgOTNmXok+HCjV1TqO06k92y2jCQQhXxr9FOGhnkG/K2KC
DIrJbg9yvC4ynGdIYFq2preFh/ihuGbiTrSwywrkr5Q+miknoKgTl/Zk+d+VkgQwhAOYnXquzQqO
13DC8QA/Rr45x1wp+SWrpWZ/IWv9fRIhjGEDSV7kfR12DZ+Td4sMVWcxsfcXmRumUdkoRo4O4usT
O53nBxNWytdjtCqDr2bOLJIKwiHOQ8xRH+rg+7ptcjQhg9ekH9F8sEQ4dbH3K/BMtL2WdOSeTg8g
9Nc8Ltf1HotaunijTJclsQjEWo1t/khy9bXhPRuRCHM2Z2H0JdLFyhvlRKL0uhZ6xwnjWUMal1lM
aNwAd1bt8FMc6X+hgFUBLrRyr/D7bRjKbzNRgW44aAVmMaD7U+M1WRlrtjj7HxcgTx1k7tliN3UI
4OJnHQkPa/b2CeX+VANmzC/Ofm/UeZNKs9ocjrYTlIAyOlfwfcHGY+/o26OIWyvgXQD67jYLau4g
5oPZdlIyBdjB5MHKIG6azG3ksA2+3d3jwR9kIzq09I+pm5mR/ijuEmLXfdDQbOu8lJFgP+3+h86s
UW0NIYJGkDtfLQ2eZNQ6cX4laOGPYESibTjspxV/ZPG2g2t2RMJYWwqxz+QxSG8xhKco/GHshmQB
xn6Fggth1kKKFzMAJEZIBXTcELhYh90ihcQFBZVq/KBJJTviR/JrTBClv7ogPA+MAtMGgbIriSqA
kLw/mtz756jP4xvqfioOkke5LijonpIMB6PRaiOmYKWh8vrD/xJ7Q1PK8pHbXroDvhXEsUkEj5cS
vbgSZNyIITfkXUqlLZCYmUd3odSNXJo7U2B8Hk41jIw2wTY7JQfbsL5DUvuEkrxr4XdTBQnUUj4S
g+RPLtWNF3buBXB3345CYe8Jmjk2JS5Y2jB9Cx7r48LPxB8IZTZ9YEpvgSwUYWZRYFb2H2j4bV+g
fQZQdqAmdoca3Z1kqkhavExz9T3DfYsGu7KGhWuRmpg/D3vekuK+W32wrvSkDYs9nZJKUvedbDKI
ngrW0fb67XrVgN+p96EpVGjClx8v9yTbiS1apUTGh92Dc/Yy+6qMjaDv9hZJNXirAYC3+6MK6vHo
OgZlcRom0s8jLhmXUqpgWe7DL0Ke7necAHG2UsXGATSqKEg6vdi/7bLAM4yXhVllnqVDhLItmjiD
n/3bFo7NvTw59fo/qGIAHhZak9Vr99bBwrNbijUWTutZIdw73p0mbd2STMeQdtTSnZ37GseI3vH9
1ozEVogBvjOMay3d+AyGnZ9zZmYxksmVmOVMwMuxXja7fj+v8framw/Y9+tXzbKxgbTUq7/ooAAS
jUB2OOUfolijSgGNcoNIF59Jxm23EUUsWRk/wTBokMDvgsLRBpW0riVW5MIS1lSmix1bpT3dZZIx
3By2XuWJ9xylp8QYjqs3k4kzCG2UJqixAWWIWguWWD6y+JveNP2GDy1ciaFBvYBfZ0QEQ3luNYLx
UaLfpUdiLuDqmkDdpOoul+4L2v2/px2cS5KUS6vCAugk9mj6sReubnySTGa50tyHNSZdITKnirWh
m/mUwrJOVYyLSkBex4CURksu9cj+91OwWFoxiur0uJq0SS1BLeYSMpT8BPUGE7iv4n3nqjBwc4Lj
rQ0bChT6E8c5L2ceGwZdCwwhXmqIK3Eq0arX3o1x/VMPBsuPMBdOC0VpCFtcrmalbdnwhZoJs6Rr
Bbn8/4iNjZOEvBb66RP9YnUCfJzRbg1CvIUroKlieNiqHJT9WLuK5tn27fty5Win10JQQio5jidW
xZSpgkayJq9jCRygzPRU9dB31ICabWR277GvDUZghv/Nw/84AusnKIqXe+lTkjnEm3FAaDxG3z6s
An29EWhruq51vlCDXze5Q7Lm6aSSVjwkPm2ReVvI9rEJCzXxO2fVdHpOZ4AB7aFgMatc/NK2b9tk
Nhyf4bPs2qsDWSb6efZm3ZD1tHt5OIxdIKOnUOprEET2vsY8iWH9xuSuS/PMBLEqzq22NRgYDJLS
Ci1GbTZT07+bEUSv0L0uNd8rGJWL6qgJ+iNY5VvnLOv0lhWaotuH+acubm05TEzVlxAPPbmLz0nT
xO136zyAvd6NABdz8APR1FDRKq+QavuVXy/REBNsuEvkG6d6RvZBkiXsd+IjMBdVFK7UsJtvv4Fw
seMPJOso500jHuvZFV5xQ9axP5hRmSzpV8Pgk/JISk4s8w64RO8ZoFlSN+QuTcNZVl5SoxIJ7Fhh
N7B8xyxYhOoCQNfiOMjzSjSmklbwD6YPaErOHncDYfD7DwF0GflzHILVkPHe8jk6b87rQXJ8QaS7
163QO5jvip+oRIdmt7G3InaF4LRoIJGWOuRMaZ4B1iC+06TfnzL8V8yfiyv2qQoZe6BsdI7DLCJL
YS+wAxn1dT2OfJWzx2QWePT+Cz4eovz6y7Y3Zb5V7JQkIGIhiVHqhyvCI3DhaDnU2ZhPuGmRoAqj
8akR1+sP2phPQYy3hmZN/dXrHPDpyTd56yd5piGn1fNSDkgXPOk46d6kco+eRaedSpeIRr5iOGIq
vMDPLQ8l5DENwGO8ANOzrs8heemqHGBvE52lReCZm2SM5WkfVByzqWfn/ikh79vM0iBGJTYFgX2B
EAiJnPHCk8x4Wak/diyLCA4srvEw52J7pK4EbPNffbDo/pzyhTiwBVKKrf/kq/jt5JsEpNAIa6um
dNzR4sW7ThPy5UApyJ1lW506qWluMBI+6ii0Ehn3pbGmm9swHeaOix782Drj899jvg3LAFCaLo0e
ilCyGCAYkbZ+ubQE7e4YPhge3Xn76NS2iCcY3xJfLWlq7jWU/+bedbFv7ns6gyDPDApl/PsPZ2c1
obob/tg6hKC8ihgDtvlyw/UaGZSS+iy/vN8jQ+exENNyDqfUKGJif6iYJ4BFOUjT6ld6I8UqyyZ0
6jPuJM7zVozsyHAniYuOjNOUYJJ0fEJnIEYc2uvKF6UOhqhLgOYGWe7cLXV0hbMcxdV331u4yYfl
MpJ+BC9ZvT9kqaUFOdQyu0sk04jcFrXvLcx/NIqS+ioUJIvlCEF/YVUCeNmsSJ/m+9Hsw8bDqKkI
VLfoUx9aZo3lWE5SBgYy5sVJX1l1mRXMSMW7zhxgkO7hfNz2x6hVRAj50sXFj4eWbjdl/rhgzWm9
0lPKIkaq9tgxEVnb2eLNVKotTnu4U1S1KGtdl4XKpj4JOI7pb/9VqQVaQc4Jn/kSUXNravNBL7tR
ZRqe8AjS2sQNmqnUg0PDE3rAYQy5FaG7WcFzfIhVjJR/Oim6HlE9r0M4RnvcehZOAnrXLHa0OGQj
3CiliN8mK5zwfgyT7AsXRv+OiIOXA2MpJKbvCnmKF7jtJSvslOh8oEPfnRh05+33WCIr6X4OW7LY
TlRdRcbd2x5OyiMnsCRFFB9UrhDC+1v22Z1/S8j/05jtI5VxYKI3Jf8sYd9d8SsauE6xJ1Wl7ymk
BOqf1SQHkE9JRTru+tsoEw5n82NvwMlwN+cEx6QKAIO1HLF1lsFxvGgg2u+uATIWgMr78O/Z8Ps/
BqjrUKkuq3lZZVzJRAz5GmsTnT86xaNhWTvjNXIUkpO17Va1cXMexs4AR/BFbZPukfTz7ofxnqOv
rzd+7pyZoVTmfq0dKgE5XCTa+pj1wLeYrL7BWE4MYDQgdvfBuyBNPAB3Om1llQRZkveFCj9JrPUc
bhvBT7bs0rni4HYywFVE4fHuyTPml+L4MgmV824oBIkuSrSiwDqwPgQBFMz85bwyylGS0aMbWZjn
zDG8xlBNgQJ2qUuhE0YGToeDohbSKkPtyNZOhj+ENekN8h/QIduaHer/w+jQTqMfEaN5Z4qeWnel
7MQXd+nY2aVVcu+SJRLyZCROKTQ1C33qc0/SIgM4/XVl3apo7JCXrwBATBEruzWODsXeK8qAlY59
tQgm+5Rj7drHTUXUkwuFXp3J7VAwNzsNglukhI0BeBS3nOPCAsJtdNhCz10EaIaorQwNPy8rRwjt
wgQ8UeW6Ha0+JqD12lwjt8OzVy6okQk4BmsmQwYrcYimJaOBF8VmArGdobQ/Q3Swlh6MfivsLU2j
XTPznr4Cx172keh2o9sY+p/RwToDdhC7Dy5uJsxUrSZkoI0PoOj2fPupKz/EGy62sDX2gjBhlr6x
8q3R9U6NNskir4BvsDuucbcS1DLe6VzdAlPw1RLN1hnWOr3iXR/sJgVFMDCHi16uJYtoabWHVlO5
ZlGn/TjjFH0QmiM5pGK/NoT5GtATh4/HgnoJl7uJxnjW1o4u3r5Y1jiB9NCtSgSufKlQJ7kTQs/A
gtANy8SSlvHbjUtkywHABcTS/GIOWpKP6wZxzBWTjtNYgdTaKd+eQimAYNkWHFMqhK5RflfYQsyi
NnBzGFawC8DzOa0S2GPzhnYylhhs1OZu4oDCdjzGks5X2J/4yvcGO6OGLWsusHvNIPsgGO+5k4Kw
S2htmUYVno/NA94aUriq9rEXsfUoH1Xz/leLNY39Q+XAZQn+J75UjIWZWZgGaQQ6gCIBiaS4g/qV
bUl6ZAXhevHBOKLWuHe6ia66R3ykBI/5zuDDDLnUHRCFUwDUGT5LXthLUnbrz9gYf+BRpj11NT1V
pCs1fvOErTjp34y8p9hc8ZOx3jIPspkml8el1IWfuDCYWqEe8phhxtUAKLCNABRIskgp8KrfhIKj
bkuB2uZiB5Xyp2c2rCqzaJHGvCcUECFBr/6u43q2ek6u7xHdIugdIDFomckRuAYwWr3PVUmHcoLc
pp6E1vc3Vl9yeMj7kWrXNN3XubVsm/aBDvZRZy5vGwzkcrJGYYchqwrfz7qyhjSRnVB2Zos2Yea7
1aF8o21pYjOIUajnJBtXAXorEWsa5MgI6m7CJ4tv1cIml9HIn+az+vFLjnXJRBpeNMKBmoSS/E9J
ilEyLV5o/FDovFdf6JnFGvuD40CYrtYzDcsFZHC3wkogCWokpG9oFhxHlfUXaQQAT9r8+6Wog1zu
2A1Yb916kqWB5VqC/wY23dknj5zc7a+09sbwWWpUlRXiOiZfMN1yYxZLnexSe0rjRA7jqNmXCQgO
Nmz45YN7PmZttgQi8rCNXkUeFtO1vSDU5FU8C3u+mNhGsJ05U7r5TnP5uNLKSYAdOPMY/qZBxWtl
hu0S0v6LEdm5ZLpgbMoJ+/hwG2VkpTPm49bySnzvYhiueGhfzK5e+SYloGMktPTc6W32e0eYr019
PpAPdByJ4Y4Mr6hqzVXQS02dirMDn0Z/4QdVealukZAfa9UK4Yje7rDSCMhOIioffliOLfID2FOz
T2dCkHNgCImeDnjHErddvrWKn/0sHXLT6uLY2+wA0SYCmTPQ3GVXxzcBzf8roCo664qiKrbSxCX6
ncH+Xm9qkmwdP7HEk0QPMgxGXF+7yeA5V0KOMsMTzSxvju6P4ctfDvd0HDlnzirhoY3CoI5oWW20
RzTPNclxeajkFnsx5WIZ2kckKwNdB0vY3rtzT/UoPxWyNrsnzVHSeVs2r5qfSM+/9WnWXwnAqUSm
IhHtlkFXNepp4hRt3TH0XruVClYA5r2/04yVpbnVZbwvKljYBtDV7hIEhjU9uZZMSt3tgOFQcsvE
4yQ49E4Ab1xM4T4+U1QoalFqI23gzYl3PW1/eBoPxtzGJp0tQ1pRV0eqjZVrfdfCzpTh9ARlqWN6
YjoOXyw75mWO3PXQAPoibosnPkL4VeVrABI0fq+mS0KHPW0mnidlF8Jg1S0JofPypOsF6Q9f5R4m
QT4sISiXx1+uByNToiTlbZ0Cd+2n2mmZOBbe/IEXNdJ1ccbE9mWOEA8n6BNUuJ6jgbZU/LasH4fp
ChtkWk38PTtzPo54bpxPjoG03ctLgtftpQY5El+xkcMxlNkifZIQLM5TWj2basegQ0HMhLlL4exh
mi+rgtV1kweaquegL2B3NmAoeMrgRLq5BmtooUpSyDrzlOcrs5mH2T1HRqVFIwiGh5rX2PR1KKdN
08QlFdGK2wiVPdbqbWMFeuL1BG3w8G7GhGXp9oMu4e7l0WEk2BFF/bG9WYn94D2QyZkpbY7bmhLd
AAzJcDFJ/88XHieHqKsN83qTT0Ha1PNF6OnnxnAOcSUlIekWpRA7zO2LC7/nFFO0r3YtP72+a+8z
kmOrKOoaiLXJzbRt4fX/1YCoY+r5tUMua+QJj+e0ovQPonhX5d3+kJFGJ0j1BzHJW0AaDVck1Gfr
G+i4bjX51D3N+RxIK9/+J4azqLQsJ78jrqPypvgLP6Os8r3xt75jMUFmtFFqCyxEfStlM0ARXro/
5SvLKvxEDnWbQDDo1pA9tsBoJHtFVN+joV8WOeFSmJSlAioiOyBq0JCDIEuV2SJ08aoz0TRALIzt
amXQpRN3v3T8LqJChsALWfDscQrVbP3DBHU5UC59cVJlF5uMhB1eaWRZvp04yxX+DVPvSMqBpnC9
fAFsHizapsN11yUf5rc3aP0QrQ/+FIeM6DteP9eSoYY9hsVj+C8oSzthb1/vVUiQwKa0k+2nhGyy
grKYNIK3koKKqKQ8o8FSo8gVeXG9wnNeU6uhKsuTQSp252NY9mMRj5A8UhtPWRVkUccgsn+0noMo
M35am+UIlgfd+MSyxf4YT/tNBMmOH7bayVZ0Uj/SU7Jxubll2Mt05XnwF5yWdVHOTIQBQwpgvfJi
nqf19QK8MxgmhcGkq8mS85yR+/OzKrCkBqaPp4X8Qjq92B4ar2M9jGyI4EQJA/XOOB+l11l56dgu
NhQTdVi78H6fluPcGUTfDMo1XKW5rsh8sjDp5G2RQgIpsz21/T/+oM5XUDvET+82KbziCl7hM6ac
qBd3qiPLoSLIYSz1yOcuDcxSwGk3E43yx4iwBlqf/vbx8KRFEuGepeiR+8ZPaM7dtAsPHN7/rHLy
zi3+N46Rb/EWXRZO0RaMZPjxuNzwUmjaKxu1HanR/o1TfnLN50rNkGRb4DTU95qyXDBQy2E816fc
z3+9l8SeN1l172CQMEoIlmYovsZrPydJamgc6D44nv4NzytdknNvMHCwW5iFAndy0/GTnpPHcmQy
OqaRlmRFg64ND3woS0qKWQWW5Qk6fCr4ZXC95oiAI1ofjDNeNr6gRzneBXNMZiScAM+oyJg4//Ac
boEN1q1BpeKF0G5jPTutJd2ApPXZYF+OeRdGSZo0N2DqzXCNVEqfO3+7X6z0aK55LmCw6rxPYy0H
P/OLSaglRWjVaohlmmwkHiGEd1+Ah4Qhqi0mscbstBttdD6B0O8lYb3WO2ekRHKI61l0rx1FqDyP
8zl2ttANgPhuqvzKLyj+R1loJLjNFsvGnfhNJ8lkU6cQwKOTrTpGlqEhpMp16WASWqQxfCReNlbN
GbG00Eb9taUv47F1Z/69GLfTLPLOKRs49YwvgJUkejCOgb1r1F3TGKgmdIh+VOmGJnc7FzP2Jwhb
eonUMdsrSDuu3+xm/MUN8eOF+qYrVimQ0uXiw0kWXSKPGpYV4VWkMD0yx9RkiKpIKctDWdwztvVY
5s/oPtt67xcxDofQ9gSGl1t+uKyXaDQliG1AEK526GtAdwGx0FigmLbyFw4j2fceFajvoATCeyN8
CwfxbZtfmuydu1rrkPJ7aKI+B5bFbCTYu2dtvBdSlZXmevUT9jlEAxJyUgniEiFvPm3UPbEpXALz
ddmLrTjR4suiNqsx2no7XUr7O4Wc6NwdFE+8KoXtBU7UkxxyfXM2jmIIcMWLzXyCCXSnTMJrAchf
gt9wQIyH7U89nqocvJg4JQbCjZCn61QOKV4rTYdXOdLXe36UmaWBQI4Gmr4xDKPe4FIvslakE0L+
FQIdWFjGCtbk6MfAxgMwU3PuKmnu+8+b7Lm3dkXVD95EZLVhIcum20C3B/zuHss9sJBHlWJKOQ6s
4mJbAf2TfqNQsYB1DVV1jzkThrKzodWlGrZ/i5y7zHcvVbECJwyQAMXpdv9YJ2sobF/HiaWp98sU
ZJnvjg7deehtq70+nbsrRM39frp6bS3SevOtk5+ewhosr8ih2t3/P+37CIS4Anepy3xn4q3kTIDk
JnYkTwO9QgQIZc+T8xm+a4Xu7sujp/yw33QpTQjcg9wrogDtnge9VLVU5m4/ve8I8r3wYu/WHGmq
S52aZ2tz+Af/+MGV8CU7oun0jkGWHYkh2hst+WKmggTOazv8/zCx6JGcwfmyo6kHQHKcO6S+xBcN
mrMVIInZGsWvIqRIIlX6803Omqutey+pZ5NsQld89F8ZFLDZWZA9y+GfVGpQL62OTkbqKVxkumVu
q/cMmHQfN0qQsiFjDnW5YpL5rhG+h7w8p0Iw4lQHDFe5e+potHFfSTyNY3S3GmqdR+XbT92XWORi
8SObGeyqZLlmSG2zCnL+6nj2jOHmNJeUWee6bH0J7j+J4vo/a6y8yuDppxlrvcts5vmRYOZpvV0H
SEgbOvDwKtkysM0zqwglUwWv2S9ujU4k/mdswgQXQEG3PBu0XisXh8CznLG/amCftpBCevUtSNWA
jqBimqD7N4TAR6hLX42MGqMvYXh5TEy1zwBGPRtstzoHks4N5EStEiyT3aYqKNb5TwxMuv+Okawv
SaeTTigeHSb94w80Ie7O4ybpPWg5SQOqTt33ko5IH4JSiZL6JJlBeuzmo84OlOJNG4kHmAooEu8u
weZ9TQ1AVE07J26saN5XyF9zr+diP8uy/OvrxzqI86zDI18R5J2o55OCQAOmhSibdO6LsmkG1WTl
x/Vr+k1diJIE3ybTQb/zh8eSgXvl0R2sz57xqRyFkn1xd5j2i5r92itjQ4MjFSCRGfdhXMFs097t
UTr/SpfVOtwgjdkVo0icFWkFnXDwikW3Yw2eeS/QsU8Qh4ByLUZE+R5+Ud0V2xoTdS/mvQdo4kOe
IgMNNZQgyRxDJHSpncdAu6fn4/a0RFivdbkN2iaj3b7JeBcpW0AZMOJKvnu2szY7qgc/rC5bNjNe
eQbGTiFjjm+Qq7D5EAM+XdCRbA9pr1XAamrH/Y7o1V+t3yfyO/CJw27gOXd6RSo5ACZh8j+GBb45
8ujKMN4ee9gkR4Hc6x8smlQgn0bdPnQTTggkmRSuSaBTjgGRqw06rGPvstKvHix9UryCoLbg66RH
bouam9R+TS6VYeXZU5QLVepteu2Mz2XDmPApLZJCiW65A7VDL7I+wVRFPSBeNzpp/TW8HWs0hTPT
DyKfvXKiu1PiDnNhGgamwkN6rXbaR703UgVl5OaWnEijYyBannXJWcf5GDG6AWkqEHJVGL1CLcmP
L4Drj0HpXz1rmw2ISPXFOFAzFHX4v4eMRTUmbGjVNlsnzEfOwJaEETIoaOeanFAVYtOsshNtFcui
fZGrpYxZBETu/xpfuz5Cv8TsuKMrIeQNRqVUVHcmxfaljsW6GSpfHD/FSIVk+9BKdDFLlnf/ZX/3
w47nabDhKZgCHZTUzPkovKMhFkr/jG0fbD3/zb/k4XvJdnX3NZcxGQiPV/etgpZOjuMnA4KUpI4y
DGU/xBUOZVE8ICWrwHwOO+NmzBoR48LZsPtaAW241BHqbJWk9AQdWiDJwO/ICPi3bnDH6l6zntsL
TJXT4Lkc9OVmnW1juBGzQLHQj1XfwbHHY3vK3xa9B/IiLYdcW00Yo9UA5EsmPvirw1NUjcKDerIw
HtD3F3wFaL+dJUEIe3ggDS0CmJUpdHegrMCrFL2wXhuqjKDxb1/71nbltjeMKG5wllBG1osPysvY
qaOilmRovKk9eNYN9bS5LADybPiVOoHcANPlYVizyvG4yUNECr7TMFoYVKkQKhfPzzN+EQp6kQOA
2DCqWFqIXo3/WQRQnipweLjL7fbHRLBAupO2xFwrjsX+vVJ6etp7FLNAIkagDV/cVgiqculPzMNn
s1taW9hNgZpgcQkIBkXJTxCY2CYCkhX4UAjTf6F36TlXK644IOS/oN6y4MvrdSSevA5ipLDnflAh
3s6o3S6MDALa/o/B9cqOmkxn/P6wY6NaQGJjOe8KQ1Ou7MwvlX+bdkoQT9dohuMmbK+uv99RyDvj
UlCIs6CnGq7m/U3ZXI3eJrTyUk+/aWAvXcaxER+eMln7LcE/0hM5c3Gqu3sWjSJSlr27uPz45TOb
+Jh5MxrH+I5koFhcwuV86aUEuzFHIHfLVsgZkpTOTq2bLEDpxTzFFQhoa3vK66TsWcFply4iR5gY
mse9VQTuG1toOiy5dlDZMymL7gUz/KbkuiQQ16RyOrvOM2ATOUvJfXzoECX+YLAhctOojRlOPE2+
PxHpR5BfzNg79lRWpexEXY3eyopD5BKuyqn0V8iYnoLWCVV8EIBQ0iuzvuNi/q+csSyn8Zfdsli/
t7S3P2R97ADH71OB0G3IRBGw+xekm0N7QWCBtx9ab6A/i9YMtEYYutBrOlC6wy0c0HvUZE4gwFLU
UDtW4l4A3ks4EvojyHY3X02uTpxGAuIgvtwwh9Ky8eCV4wYfTgjvyM+D7tq/3eeRK5fl4w6zs5dK
+9Vojt6382GTE6SEpMerauFrULm+/XA2z3Yiz8AHg83P9/c0Z+gVfAyOoHUAEB3s16I82J0//rth
C7iJ1oKHtvDABNw/tStWpeX8aJt2OYKFCNr5gJaeCKDseqO9FwIOdN4LsEMW4EnGm6CYmZVoSCsv
qeStdpmpWplp8V3qk9zcqMRvXRIPdAunJHNwvJuFfyDhCPP7iY2dSR/r2esKQiCeL/+gSqAfejK4
i5uuAi+NComWnjcbqOYoTCy/Dujd61pf3ObiHQQBCNlJH2ji9mhQ7x6NpZcazO4zncRHY74kiEFm
9VBGAZgDaGpiXfnTuYbwmObCiKa8M38eeQ1AMq0sK5P8ymfuBwP3qUlPLYhphLTTZ6PNTat6HEez
srGoSmuSENpSvmPkWemp7r8FCQsb3tKPWVw29PrgzDNQsvQaeKcapfo7c1TAqWURBW69Xkg//A6V
gpaiz/V6GQGyaGsTgahi1+sNY7/s1GvyfAXqZangMV7Z+88/GYadefU1RbfG4JgTbNxRehMdUS/h
POZDF/XwBdW06dh6Ap1xbl4vG9T8ZsHtzRq/c5MEvtcrNkxMq7qwXDFA662HlkhN4m6C90X46NTJ
ArQ8rl38HBF8pZB0x1Y0fjQMvIaEbfch8d2Wb6VkM6r7ZhupklrOEy+84TbNkKwoRpdTyVDhOJdf
wvO+wM4V1AGGQMtlAxJH7DPqFUD2V+FdfnF/AQdHFbYFZrFWKSkESPSbYSASVgdxhyTG7FNDEXSd
bE3ciujgQvv+SjqBrIMfBm759p5sfztSnPHGKd72OCERIqa8KDHlRLRSAVWsAvjTMm/dpQjYR9Ex
j6YGnckalBftr9OmgvDKQ0Gor7AJHKlL3n7FqG76QFvnV/KaSjKxlrjiEi6icZXETKhOaq87e5+j
zEgWATvFbp5MWcZdSfg/rAas+RqCMtYgfjyy5vS4WkpO1sFt16eUbHAx5rC3hZhKSrzYdAnwoLIN
XiZJynn30uOrZfjgnoNrs++0KzST4g//WLh76M2SFmDqeTe8wf0l4qTX5rWpDRniDCaB9Hi3fSkR
ZEh+ShjuPhZ4BenoTujI/HS6BbBK0btA0mxAVQdZZaA/vaenrUyA7GP94+yAi1z+E9mQbED0665N
oThtfc4iZBOARPHqNXhiMD188UpNgzO4Q9oWBWn0DAQbM4gRDI7A2QcYMc7A8v8GH1fEdyi/WENi
7i8HGyOrn5NzZ2s/SXNuIFskoj2qQk5pfg5GH6xJFLvI9bmv8BfeS+N23DDxExXzOSkQOIiP9kIu
vAeQtZmiWqmyQEMPIfauphARwOC3P5QjU+RG/aEIQMe1HzKoSmbhgLiJS64K145zKGsK/dTy7LGD
Gy3TpO75mVKo3487idrXQ6o9pkzJIwlcQS6MxdC48zsT+sxhi/YNinOnap/fQ00hHDVZ5CmCrTcv
KNnrLfaonMq12JMeWvsnj6RDiwURfNShUzzAn37/DEz2jXviVcg6xBHHZ8AaclvqNNNDyem+rF7h
mWp2bk4vrJVpEyrMzDq/vVIYs6YPHEjbXAJ+9Q+3j9u4HiIStUkYCXyu21zu3rZhrrwPW5DI24Zs
ShNpzdSf02pfjn98JwO+7Y5svqkMHdl+jNCbQP0BaCzB8UH50kHXXFOYZEvl+Vdg+op4KzpTyqjf
zhE7BwTRZxJ4d2kwOwmywykdvGg4rarCblsHmG8TyLy49QsJEzcyLX4PWHQyjI7sL4cMAjiJ3P2W
QMKnX6fzbVxKszq3m683Lg7t7zIHieEYOfB8vPb36O9QcYMIKNXd9SC7TFQye6iG6dkAyXNrk5fi
DM/JwsgdF533jJdEDmd10bLXcLUftkW42kqQuwhRyuXgjPWSVddY89C5YCvhz9fQKwPsKtE6B6dW
AlgAKAUDj/GXQF/ulJK5w2oZIkSE7nEv1X5X1oWRWoVbiz17pdTj+DF1wICJ29Niak3u3Qc8LbBs
Ry8+vO2QCmVPKGH0bnEggjIoD647PnmyVJKOTUy/BcpxtubZWXona6FMW9yOPnxLXsGpYWAadQMa
7pn/UdXmju/GMrvB1kQ1IT7BHTZtCh5CxmUMvc27k+MDkMoOdwnI68XM8qCO2dxv3s1RyFNLr3wx
86o5+2wSieMsNgODOapLqdhocmWORjpVlPvDF1reY+QtEUiAY4vdhuDvAdK7OEcYeipnECrU8BR/
VY9z6p2mODtzOS33LpOKjQ67Q2rwwH5LFRGkhMG1ptagxpEj31gV0wUnx5UU4NjmFSc9v20w7fwV
y/yX0dmamyiKI173QvMQE4n4miYu0cBJx8vFbuubHEwHR2xZ75CIylA5RbKW0UgdBlcOLDmDqkTb
on1G2FKquZIwbYNcgdzycTwvUIV//RqdsSmRm012kkZ+4hkIHzwqegauXNOxoNblPYIFyTVA+ow1
dlESAN00kEeJNweWToTZpiOjFR7MCduSiiPKvz92roqpuIlYEriQY0I9K++yk4qksQ2D26utLpUc
bWzEXPNvtz3aLkwrm6l2syEyr6pqHjgHPBuOpz9W+gNdhs15e3l3lmL4lMTI4IrNigm0YQSAW1gd
6KRpWMX4o8ohtBeq6B9BPLUrSZ3nBSx57NPeI/AQIeZbx9NQXCxO7SG8jQ6p5ifYEahvCPEjy6QA
bqY/dXYslj4OXs4KO0l8m2f0oQvwYlKqruXCaD8mgNLKwRQEGGduT7GGqv2ojklOKZev+zaMyqWm
7g5JqfvbJ/zLHRV0wF/o4x4z5GJwWYTA94ZdKswwgXhxBxKShN1R2pKQunAm8cfC9YxJSQnkBsVs
YfrzqiL9ytDd7d3zfG1nFvy7Qp78F/mSctvTAWi1pMryqnJw/yoUUC/vSjv9AKyaBskAi7vDooPI
so4RNehIyTNbKf024yGgfCCKJtwgXgUYhh3ZOKl8qxxh/dx/GccPIVVIN33TYBJQD3HmXTw8H0r+
yH6E/K00VD7iJiIbl1PnK3zmLY3vqJUyRN6Mb8e0GKSVYQ2gir8okfOd9rPa+rYTsw0Z665bqBBm
gKgflMRyf4Tk2ffh+w0+HyLB/SJ6qAF6LyeFIRTFB/FqUfNVXxOpqjoI26+6GVfUXl2TEKfXZAE8
VYnFPQPWimt9mCLHAu05Ppyx8/5mnmKtDU8dPuCuaX79mD9jVbVpnb2Vv50pazJdkBt89GLH54l3
n7Y4KTBD25YLbr1O7Ttp0jNM0GoxiDyLI60WoULw/VXtPGX/YkegtbFKyASiUy/j1cy8VbOYwlnR
M1q/1tmnvZj52+Xw9kO78Q+fi3imUJgQXd9ovFdibtdLkMdaIYeGgyJ0rOPthlrVpnMihQcoXfmh
l0fLkBHzmhWLOVrv2ZHC4ptJUUFT0rKXc8lPWIXRQn5BfuIXTHHx74pvYelbAhtOuv7WMcLaSgeE
iHNKzRsqf4B4VkQsDqadrCYxlxrU1O+9Vsr60vusbetGaZyUfXNHTVuGFKg5GTa5sk+ECYJr5FpF
04g9CfdktmlF1vVDBWWz/wLtgQebfb4nu/VfgpBNJtVz2DIV0IDy8iumlj1xWN7THVlDprzjv1Ag
cCGvJsPm+/BVIX1SuKqI+xaHNvud2H5/+AXlLBmrClbFRgZFjHNuoY4q1IvfWRb4qKhB3ANUCkgn
EXOKBdGG1XjubUQE3EdgvULaCgyD71RV0o3TRUdHoVkRSki9UY0hrClKF3g4Ik9+Tq+S8QlTxZmi
8MkAbnBFGS1yEFHmIVpoMZGA2Smg6K8uS8P/FDlwyL9OrgvpenKPcP8hVM3CQRbOUvT97C/EX0Kl
jHfZFntHVzYESlyoByxQmIYOkINlCGpfQT1ek4uR9IHVWXzVRSEeuycWGcASRnbYrBq7YQWkIZUm
nR/Fo6TwnaIAGG+AxdxOqzBQiu+GEJfYtkCPlY0kTew6rjYYAhhY6l8YVN0uRkpSGddagIVPeorb
iiqU+2cvygwvpvOdQs1FlRL7QMJvk5NTGNPhTXJsVXgdFjiYyQksVz36d2Qy5EP5KhFytzQBMPX6
og5gk5aZvqboZiMPyTHY8Dl5IvL1kt9inklDFGypWHSeP3AQXM//Adp+L7FMPneU7rcOeUtIjn5c
1gcT+sPbxj04Aooue0ZXKLf8U1AH3gVVuXUV1hoWvTGx6ZB9CGgaspb+CCC9gGaT+Z0SebrR6pvB
WlEy9PNjjsywXCgAEXD+nkkcnXgaE6WOF4kBDOdRkc7Pm7hCg934HvKevv3mEmwBJFv8q2jL1yhJ
qxwoIL5hlJo2VIobwBhjlXt1MIDDDCJLH+pW6m0NYvUh2u9TciGn9pcvwbP7YPUT9k7bVtr7SJER
rvjiQhjbyCxkF5fQQa7qPpQ4pXdtQ+I8OYIsm3zrfrwEAdmTC4+yEYoD2jIRTmPP5QuvLgPJPeBt
cmjlGeMuyWADM6V9CKjhflo+5Rf5vGEqYQA5PVmC2u0YLmPakMTRqBGDi3kgohEtWsNpC1ujFc6J
WE3y3V8y+si+lxyrKwROsWYvyAWhrzdCqYodt2OtJAPPBCvwWTtYaD38CCr//rQiAgzXVBLEyGto
Rml2ppfrxDLji6cuX2XZINxg1Whusb1RcxpJMp2FGB0b8fQCpuauvZ9/vWSHg/MlbHGB0RCi9uIf
K/MUcPURBA+Gvzprk1l3YxwVBdXyiKzg6cvAUc/T+vkgrdgeDMD8TIVn2qQBbcmejt5RNd7DNbRq
iu2CaYcvJi07XfArQ81lev8MS6nPxRvnO2XwdVpkP9EJeyiGsGCSiYVaFrzSIHk8Wrq9cDFKUIEo
ZQAib4IAUEHGqMJpBbSI1Aqoaz5PQWg/NK6Celzzq20NujKZUBsoYyvxOWiPpNb33aCWT/7yMd94
/VK0w1Pu9yv0BoA9FgXz3ZhxEVLs/YDr92OGQZb8pvxpvuiQ63K1Fv4G/GLss8B5PuysZ4+vSDUw
FQXPZ4Odzxh1q+b34Q9H/sKsVyR8jjcyCWgyBGAkVxMyaGrzzCGRHxDjrN4vNH74xJwImB/KhtCw
S0ORuIVP1b+bRyG1ohuLh6JeT80wYn0u+bL/r7lGGrpvHakScsUJcRowl2V3LZMmVu3O/Tub5D4z
h9FxtFPI1HycmzjktyBlXgaUwAQDSe+jqGTQHNCwcdqPFDbhGm0pmXjqV4nf49PAFV5HvlIkLT9T
jbs67bdN7FSefuomG8XgslVXVZT7LJ5Ei3KxLmrlIQju/XpaGwUgDBYMc4wVYdM3/ZhF3UzVzbiF
CXzNmMDdR+X14cuj0HuOFOcyPCKt54gRVHdmCWVPmWY2gVGstI2fHouJjZKr5YNOepZkNbBV+hvF
ZA6u6OvwFAJmpidErzacLMyDFSkRx9sJ6laDDAE1NR0JJwsUL6QrEEVuY4ANhniY8Sv2avDuQLl6
kzkyPdLnF59axF39vCKVIfkgmmw6P63F0fTbDIjmKethbBsMm1e9GkQUdrGfsF3DuGN+a60QR3xE
Kcoe4pq88kP6m0/oU4BadGv4rxUh/Kxm8ZRr2Cfei5soyGIs8jjJZERTyR4C1zwCjjeOscTgwg3w
66WC5s4L4z/EbpsHS+qig0K3RXIkok3f1DzbFIuC9zkV+K9DrJtSKeQNcgR0fsAk1FcWxKly/W7x
qh0J6uh27u13UxtLjKF0arDNcRQyKsQF1f2qIU4EY5iQUIpb98X25mMeWlnlodYoN+Gl5vKfp7wr
XYbQeRtK15VgahEpxKOG8usNnBrJkyd3Mgxc4R1DK01kPi5OwgqoBFKrgUTkFdk0zcS5JHf1KuG3
DgMa4FsLmib0guAvwPvQhpUlzigPgX2TJ3t7XgnGa5TwE4hQw0PHKTsE38uxh/o5gArLqqXc7Nho
C+b6l+uROX+VFPZABzYHzPe7uxKd0mKUCtKDG2GhStncBVyXosREvH0X0Hr7yaPQTN6DtOYIm3KD
lfbOs+pfKRhnlfbKSBEs3lADnbfSd/XXED10OZvcJ/0HLriineWJycDgHrBC1aq1iF7JWjuZklrH
g1HBmg+cWA5qNE2S7C2b7yu+CQwmQxjfXusrZBuYMOaJjAd+xFX30/B8guM098gzUgcI6NIemu4N
cKr/v92sTyY3HDmNqXuPFc6SfP2Fu1JrtYJPDhs4Mp2jY8LKdkZzjIOQIz9tAVRaryvvWcTHqfbb
hRZ/g7cmfWZY9eKXAbcGUbFSM5QSkVSsNSSVJL1vDdYM+iygKT1EZBvqWgzvOBwR2b8/geiFZBar
xcYcX5OCjrxqW2+Hc6mSaVaRA3f1WwT8UJaGsgAFg6VNbkclYGXMNDqWZS44UehvXFMPauZKQmnl
YKFkeihymqilqzb5LpzFT1cp2rSt8BG2TR1J2/yYabPXzIVqgR8bez4fU5n3PN/Utg7gPXQaXeoc
zP1vvsRY2nbjRjjPdPTXam7w/wcclDR+F2aOokJObpCnR/D6fVZjNj/FfZ/phVqYZk0Qvyt9M6eW
39osJ/mjjp195hdDHUBb0zrJlK+Dq7A68M+LqRcpB/9jxQLQlGY7M3jMqIFd+LRy25lbOJIdwARP
PWT1GWzuX5rfGJVUJ4A3a4THe56B4jKKL9I773JGNw/XTeTjPT7xES5Y+lHqB6WbCeSKeovcPT+p
+evYcV5wkdIVvaMNRS8ToRbkqOI5WDF7B4nAhi0pNzj+siWA2bXdJckJrjyAoesPLP//mg0+OMzq
1mqzCGHLqqolvLsVTd+Yses/6gt24p2lDp/4XmoonZMbsR0qB5eyRQCuirq+iE6ANz/HFyKPur+U
pPkCfx6oaBmx/Rwet5ieuaBVULzs+VSQDFPPAOScoU1Xz8uozORoera3BqIjNBCzW4akdQ+GNUok
T3m4xdR5U0bcvKIzhQHZgOzBupfgh8iPzjdYCogPxLFPVK2eixUpkM9LKM8GuAxqX+j/l+TxkJzI
iV6y7pqs2O5gaCpBHIqMC9zc6+LqSFBHCSvD6k9Y3lT5zNo4LYF9mFstHWdMqyu0IOXfcJlYB69g
q8QRyWmw72w/wZ33+/zdTzs1wMjexdM7aPsUCPmJ4A56rx69C6lKiP2iB0oL6ouzUk6kvu/e52+2
6sajqOX/5xzLSxuc1wlviKvgHETcO0f2a1RAXyuDGllEVH/olzXrsbyiWSByDYKujoYrrIgyDhDW
2sUHOFCN6xl4Y1uL0SzVlB2IsyRfSCxkCskWNYZSi0puE/wOiMo85gaIVKBsbRoeszPBC2PCKPAU
FcXjlHlIPzcJ2ac6U0PbDfp/DevsL7NQMlkXlIUSJGXSAedfdHeo8+AMsjiVCA3GKNQ2JrJ1UEoa
rf1+AXiyoIguJsz/EwGCIDf3oW+vM+ecrAeKgPEmVI3tlRm8q4RweuDfjceCD0xsF5kknSgagI/k
lLZG7f60OyDfa8xEQSPGT4gG+WSZf1zcE4eRqVavMU4dqSxxbKYGbOLafXlnxO6NMAVs6TTT9gqQ
fSTKnrcyR1NicVo9wpKFUOWHyZncDFXiLOeEskKw/JsHYt+kPJonSH0LQ4y1vHYGWRId1O4oM7It
M78ZXcZZu/uocHSX8FUYF6vOPCtCa0dE/v2Lc/oNjJhzkiO2iMDifigRjaGvT2e6KGnCkUPXTyyM
xlQ7Q9Fl4DA9fx/lnHmCjiosrLi/EFz0l82/eSq4rQd6LuR0WLYHvWta+VdpYgNwLMmTBYgioMt8
wJ5fA6NTnwdlPyZpwZkRVViuV15EgSNPf7E4vDklxAFo4Zf+Ht2pbNjhPfQtqw5yHj7CrNF6lYN5
erDRt1xdHG80Gy109ZcNpJj4Qfy43wrlnodhGBMeOzTCwL++WV0bibtJNbaMqum2CfNxFSiNBIS3
lOxC6hyA0qGyVOQZ1SdR1qdH9qEYuSDU5Uogmh6w1OK45KA4xo9ztTJsS39vT9a7DRCz+z1bQ70c
fAWW0h6ZbRXs5eDiizenquUKtjhFi4Dj5umsw63HAxZKPKGSbMNv3xzehsvZcEESnKlpi1PUENwJ
zw6jIpKtYSzr1zSzTcxtLjIQ7zyKu/eQsza1X0JJddeLik1Lr+zvKHq8I8M3hNKL20rbQBY/emwK
ZKYQ5MRRliirjifyDYkCr0pz6JcU1FNDqTh37gz9xF31bGBUzRCDUAmx8qlAL4iJBBVsfeEKuYwd
H4wnxRIEY2Fv5glnK2sr0UWSjuDqVZMNhIYhsbyljFdz70USutf34yAsZa8XR2DlDNmcrocFI33F
WbJW+S3bttGBkl65cq/31aVibWD4cp20zPLI49qFuNygCRv2rzgEluf9aO6bMhb/PrmFN0x7YL5m
cMt2j/KWzNkYRhd3W4oGniRhAT7e/qMSlxLnVpfwQ8J48b+a3G0qrGz4tUdb/CDjlee/PWK+KgsH
LI+g7n7Rcii7KSyHCH1s0Fa8tizPF6Jiau8deYblWpjfsGTyEm8z4VGpzor43F7LcWjchtq9j0ZB
K/jslDzlq02CueYxt4VwKIQO/E1eesLnl1cR5FYBOq8Bv+mV9RAkRUClD+dD1z2TiH8ebFe2eD22
L4E9T2U8tDfDJY2s9mmz++rnJ4JQiOE5uJ8UZ1qqkYKDg6hJFOXsF3GspVUWskxjwCW2FMrqjaS2
a5rMLsSQIH2kv0k3r74DPYJfCINYpcMH2+wxeghixSyXvRqieA2VHdHrfUa+rqpEyf50D/lzuHoH
YWpIbXZ3TLVLftYR6hJMOcKSjIyUcUumRXHhT5tFZvyx1N9zuELOh2Bey/InLlWGXBGIXLpLszt2
tPZgqVPkmbh7a4jwDo5ONbwXYRzJHFsKdjN0oMrlRMWb35SdxuEJftsnPJuvwf8W3l72qhihdW0B
tT9/+GhStO5dl8Nr+tmZAfG+bjzl0+EnOQliOO/KXmVUnQmYCMRVJeBZFfZ4x3CUweK1h4wWGDiI
ybtnMxpQLKwUaufNcoPRsbvIbYHXjY7GIoEhiLYq2qzEyQzpq/9wu6/q+kpfDFgIeRdDfHvTkw8t
Ztc1M/duPwk7oMgamMD+OnKGEYNhmxl6DBeaZb1Szx/uKyNcR7bhHHFTffnay5QvA/EQAK6XtO2j
4LmJcfsdSjThDfOur/AzzbIxCpXM9WjM6uPsCjchul/dQpnZpyhj7j0cmfIVOwBea5uwXg3So1Cr
RRjofSlT4cvkhHHLhSLJj7oKYOtCCXQSwKHKRPLFNHOrIqMQXxQoW2JzoynAwW0+cwpmJwE50PVY
ImoZwiiVx3boFU9tsyMNTwb5jsAWngWonRI+Dcp3OCnZX+v+aZf69WFrXXOSAgJytDELSzFIoQAr
fHdkHPzdCLS+0S/PQitp8E7YzC42bwFTHfZ+qy8Lh5FOaA4mZKeHeQ5oJv5tiqxgz5ET8vAezK5O
ZX0fL/hJOS2ykk/b/l+vJUsSoXKqNQw/ZC2qwzedpncQnxox4pmz0hM7kAIyLt0yBV0LbsKeWYbL
oFHnR/vIjKS3OMEWKWcKDrRm9ChOFiRY5RNr8cC76et2Zd5so0X3oNWsWj6hU4ZHf8G7nxJ/a0FW
Uqd0KrHpNiElmJ9P9DkUU0LBLiEkDDCn0rvHrI02Nas5/SypxLhwPZeE3dhFLC5x4tXLBlTLWrxw
plSxKrPuEifRJAVzZ2wfqylUEAuEYTDZ9+snSdDVwXm1ow+x8zavBM4fd3bfpH27uwec2qPV0x2k
39jTVQPUkYXmNuM12RpodNr3TxsZo8yt7uy2X+uSDnUXSHwjB6zeQk89ZsZ3WA9Xux2xWUv9CFvg
C/o6eTu0V/SfR8jG0VvEYdetHQ/Lr4X5g18P0YrkGkDsILHUa+d9cTl4Obq4A/pm2XsSx11tiT7y
IvUnce8xba/kH78m+QpgMXghTxET21y2aPFFh2YMxzorFKuSDlDvMaOshHsj9h1T3LzmxEXUv2RL
Bj0xuofmx+Zq7Jzf6mkaHdh4OvuB0+eKpvZVcywW/L0Bw5O57i7pc9E1+8++Ug8mD35FPKvhZA86
kXqAeOvz22WJdGkCoJiEf8ypXdtc8Xm9wXL5EFRuLmQgU4X+dG1OEuV+PbF96WmdJ+so+GcBiRHd
T6VaDj/9878+oAL52dVM97cJ5aN2V4C3LfpFxlJ5UuulCZBY4hJJrVzR3XVreliulT+ZoToslNd7
QQsyQaWkYp6iivAIS2UjcXIXXVBCz1e8eXDhSHtXl7CbsYmXdbRmn/xGm49td2vrOX2Ufhze1es9
r3qo0xfTleFcwM4vYtoHDWciD7St0V3LM0z5xRBz80ikhM7jBW7J6uBxqqFspMKdZTFo1asZAYcJ
WP2XNI0BqN0bYpXw7ev2l/OzMq6/ZvEQR/cFXijLNkzRE8zXn8JVqZ5GV4XjY3fVVKwL8YcR51D3
8kXNL6KWZu1OBGyxS0ZFwmE6k5OYv6dBS5o2SE86whEFPTXb1YjqIPknfWLKHJ2CvWjOJ3fDPOmD
/HIHLmol0h/ntZb6J9wvDG1xY82nee6H+CzklJR9WTOYRF7ZXZU+a/je2hlkqDRq5uC2LibDxHDb
GQacozqhIP3WVxbkW/XzolZ3atoG82dqmiY3Du5eFOJBJN4x6+qfi4azjElJM5bnbXwxyRudjknV
eudY3roJeSNoaI2XUmHgw+dVYc10WLRAncN53yUxp2D+nCc42VSpncJncMeuw8UcyxNdg46fz1uJ
aQ9P6urOKss9mds/hZyW1yeoOpN0dZbUvPbumU+uGbasNI90uR5vQjH49aPCvE2ErA33kAcPdA9a
wpaMJjiTd1MsJe6PHVZIu+x++ry5vcJLku084ocLxEH3j+g3WlQC+RxSdgd3gtw5eKXBpbhsTsQ8
HWAXJaM+g1qFkihwp8beBzbf3+pAL6ZQhZuSPXh0M0xq66v4zSYC9uS5JtIrLttUTLONh+5IJoDI
T5cfs4rbY/kv3eWLtRzGztQUqKd6ADJZpUYwzgwbpJW290uFCIpaUuSYZZmYQmcBcEo6+i9QFR2H
rEIsuGyf3ZKR91ggcqcSoIgzZCc7JL72LLcuuCbMeBUkbAETYdDrzuE0miQb6zYfYOt+RII+sIPH
FmolO931jLp5ZAUOuD71XOssbKRreyymFvCAzOrAwv88XJh76upf0J8w2aUbxuh6jz2XKb1Jq4p+
q1vRhvFA3gWzeTE9WjrM5hsHv1fSJZOfwfEfb9IvPPH4uLJ+ZGj0zwgI0tYMFhhKxB1MCKnfKEdq
TBbEdvJVqpQ62NzsqclRr8YK7W35Jkshc6MmJAaR20yZcZgqFCK89Od8rfCEUtxca/6phQ3jfeD8
uImth6+JJn2bK34o7mbjMidexcfNTTMdNe8OvvCn5MRwziOXlRjlmRhANl/85SBy9kFB4MSUwQTp
wMltxoPavksbOf2zEqBXEoElqm1LF5RWlwkk4hkipVCl8TKdT95Fj9i4PpAL1GVi8D2N+Wv2EY/D
AXYUKB7G2LbaI6vz6NrQfBrOEBXtTve23qglJfsqKD1gp5tBcPQemuZCBh4dVeF7VB4YWSpe2waP
achQThionpvf33RpQBXntdIiJL17CUtefe6LeYe3aSf1RrncAUaMqHgEDqHx8eU/2yJHP+dMRNHj
PFLbJafqUSslVKw0ZV3ashml3Ii0wiamcEH0ppGAdv3E6CXeOjKEBJ4Fyh5N+aS2r30C5VNcSfBk
OeoPJHUpcBJqgeqp9tU7HyBBN2Jv/W9fvzkmEPJIdBju7Ln+w4L8C0pbHZR5/Key32/dOGZ39R7J
rKk/9iSbzK3xltBjvBzVa1eAuIklVxlGV8a+iZnraAftFaRHQzl7nxZFZKG0/ubLkA7wDB0hmMM2
+PKfq+MEgJfSzkS4t70SMlT3d85jwJLmHURB0kmVf4TxFZpksVMy3gAfC7A51kZmD4YUUeNc7+Uc
LCOjNcmqYLRyvDbbn7K3KGgMzZrRSO2kNjhX6xlVd+sHkeLl2W/u1ZnmD1Zw5+CIKrku+XiktNpF
2Zc3IsEcqjVyoY+j1PQYWwIYULsu6h6G7nwbMRAGttvusUmOqmDEr4l9DTgW2BfcN1mSCkrhg4I9
C9ehxv8oY52aWveTU+n7IJcjaLfyjzOThmcH1pnJX0aMf0fyFVxBN9tHkGmDJzVrJPPiEUdlhYIY
MisJaNHdPl/rUF+HVeoSrhK48S+HJM/T7YcaxONDRVjzd6g0VkMi1yEDQxciNwL0wDWV8GIX5d07
msfI6BRiXJuyoR8980Iw1c4A7x9JCXHlKSaYn57gkg4Nw0UO1q4gRw4ziGpcIDwpJIZ43a+MJI/J
BF8AeAnV/jReCYekyDmyMwmk1qzCUNSy9/wZJ7/rdY4IuxLPRqgSde2/J8WeoRy8nsdYLTNpFQgV
orUbO5/PhamRa2Qa69TLTiKbjcmytS0Yg6xdWdqG1Mt4gmgRwdoPdFwcxRWgKLcFbWoRQAh1zsq5
AdBg5m9gvZyJjbxKVq3jjd4isLO+HQbaQViITHftzggQDj54Y1VvKm/VqV5r1rfFIz0yzLoEHsd+
iHChusNwJtNyjawEIWyoIrqoEIOL+lU9R5e2ie8toVm4ZjqcoVMalM1fbQuYGSHaUR9ZvlNGmdFm
QPab7B3fV36vBZVfNeVbTMnKEc9VoJTlUuKOXeq5w/A4B+KuKgGtZX6v+DWWnGBLboUtvAlo+ZnP
QwIHMmgvg1m9LhcoV6Fxh3j+lHiZcR2W6ePMhFWbXvifuDvfZ62YPYxK+JZMEnqHuo1Rmdg1cxfT
ekqjZZJT4ofToF7+2HHdCbUgoTMhceVEq+GFZFf4Ie3XBcFo96RwJAN0aJ+bci0eEw1d6ZUW1SmL
DRt50tWSDDGoOW7h7tq+Q8EjVvA1cD1QBoD0F87Yu89lfa+HOu48ueu3vCuQzV+GcQoo3sZfhxUQ
lWkRJmBQ/uiD6klg/MUc9OPaoqyR9WhqLtJifYite9L5hgsw5b3sXwH/I6kI/BpDQa50AoznRdlZ
OeIZMsg96AB/A15vHKgxhL9eNORAGEBfjTsaI6ZC5xY86WexLlq51G0eAbk/5hPPEd8t28tk5HnN
p4n5nSrye8d6FnKuPLJlwPZ/6ssPCZ4RFRJrZPRP9cbGdCzotuG/hR74/6WTEN8oPVVFBFJR9CUi
O46dDrboMQa5ZMAk2DP8dDArTegt8aWg8KP8Gr/VEfFVxF8DELk7S7Sm2s4z5cGFCv8PHffg0giT
LQOxSNnZjrzHk4H6Vxz30vgrd2SkGdf1st2dDC/z8Vr8cpYDD1zFVSFvriq+taCvbcgYYcEy5nF/
Z3IyfJMDj9PF7XkD0jL6dsTsMISwNM4Tu8B1z83XdkBFVSFqeRScw/LOPIfmSiEjIMJYt3Aj47UP
oj6oa11ChbKpOPBizdbPZFUO28ldiYXedcf7zUcofeHiw3xn+9w08B+xs7K+IBVM47olq4GuZSAT
ytTdBFWwAUDgFZNtH3Y0ehCv2WiMToZhkyb76F7QbBsapyR93BpfP9Tx1Z9s4MxCGkDDrio/d6E0
gElscyzVkBQCZmS3mPkEzyqp0guhqFdZT2ski3YoxwaN8gOhgMCSx3cxAqB43Rf4eqj55i7fM9Q7
oS4yx4KNJSW5I02EIciSgoghRmhvi3sys1PkFiEvBrpqTq81GTJgMWZ77SlzXGZCHJkZ3T3Ps+3P
a+/3e8cIGNBVDnFtQk+8fU7x6jFRARi/JRyG/TyBws+TV0aMrmyGlSxJjtgjrOfpUi3ddmtcmoCG
AAPR9kndW/YswbEaVD1QHnyzY6fgGd/y4PfKu3plf+VIJHmzPjkHd+OvPeb2RtrrYFCLXmyf0wdW
JS53wVirOlmGGfCrYLV4TS93G/xU64XutvnQpcZ1zXqTkilmlvhFVE3GhdA3U/BWChu1A1zcrrph
EbJUZmZ5vi2EuLOqZyJ8KYxY1MR2dmcs9G93VUWmSk8lmGmgXzMS7rHNDxqaHErfsY9uM3YlVkS4
LvcytLz8F5gGLmjuaPM4P+dfJdzIVoZ/XkOyO78NsvotocusaEIhvJIIShnr8KaklOpp3XJ+VbN5
I4tHNwW35P2ebBrEEBaYy/GtjjXx78COGV6Jf4r+s0ITPGVXLdLlT+smEvN2i7yN+YFQU5HjL69t
TFKPD51/9FnnyIc0jLwX7lkLZFJvpZFC2tgsE8pE3HMtgGy7XLMhzbqbIX9ZwGyTe4pQ1jf5ykHZ
Tpg8Pxy+dh+wG/2by5k9gREK8KDVNdgHRY8mmy1x4HlNhJ69HRChhkixZ0FDRxtAQfkXAPb2KP2k
D51WSU/lJcIckiZMj1CjfonuddSGtdooL3iV65w7ym3XHuVG5obWAtM8AmYfiaPs7H8cgp5MN3M0
iN0QewtgcVz1MkNbLgQSC3NDCK7tNnPQflJLmlujWDJMS743iNmVU1xJU7t4grY3Zg2ye0wqwseC
dXczqJJL1GehAfscFYh0WuZE4+sCX8LUd/4jJG1/eTlKzEvwNcWywffEyQOwiQTIk/eIW9bS2aSi
EP2wXpDs12XoSyLfC4xdCghvDxmhi5lmwRuwGavL230R3PF1M2VSd0zGr0avmvk1iLVw+MDBK+P8
YBc1QZX/WiJkWrS4+a77pW3qc29ou0a1YqAFOxtvKsY5j+3k/8mm/I3nycusPpUQqdncuTHF+sMj
PKqsCYcrpGpGFxoQOjFHzmccjnkDvDLv7I7AndCvBzON6W8kqIWe6kPW313MmYL8BVuDGLPcDdkb
W2ed6FlYaI3JfQb2DsBPya8qZXdUrHIwBwbO4in1Lqcb3zuZSH2kt0TfuKkwv2WhBZjto0ZJR9yN
C/vlakeQq7PcebFxod/VJRcvlUtcz5A9Y005SQT2VzcbiGsN16V0s+hMRv5J2XTRPCz9IvNEh959
a15SaLPZxr/KrtOLkxCEv2vCPyKIRPI9/pMxXzUAA2ASZAzrS+SLoUl3Tt0nD+CNGNdM8IssgyXh
YzMzB3J3cZEJfAg+AeOH/bG+rSMazLBf9blcYMdNSPMN09EPlj2+IN3ZKjZJ+8WyXnfxk9Eb2jKr
Pa5zv0Fmi5Zubp0kW5IA28YK0VjXcVnEFr+JVPT+w2LfNC3CniQXsH2r+9qPl+cKddaIwc/8F3tL
f9R65hrZIGk1ZXAUsUINeCFUYZqd0s8scBhhbJj1dSrfQ6rbkFy1Xybzbr2NIJ//WG3IJnac8Hqs
WyWq4ew1LTCEIaR3Mk0KdXK1hzbQhUk2ZXwM0GSpPT3/HFBdoYxAgmBbDkVAI6Q7dDnpuTy6a8xL
KGlt72ddqiQoy1nhVPtIJK4GFAthr7+p+GSksR1fDrrY8vT13IbHvH1qKH8jg7NvH1Z+68/woKe9
gZDb4j6vHo5tlZMKrJm7nNuGDq6lTzu1hcUTSxE+bb5LJzBg23r3W61i90podDt4igPjOGcpAoyv
VmHB7qFcTYv76wWv41k5GUD8YK/RzkgxMiw/bA4GhSofqFpmdqmcWLUgrZy/29QpvPR21nyB1qVC
nt8VTfgePQOh7Wkvrp839GwC03xqCjIeVRTSXhXzXyBI2srm/Uo8eXA8v7ko99YTWRPac0WQgqjv
3Szb2Adxl3jNlqApXrbJYSgDu5EBk+dEqfG9eTSx1De5CeTa7gQffrEXsJf3ZJxvFIsQXew6oifx
VZ0+4UGO2CPd7Gjk5nhBG90Add9lq6jBbX9837UGiQ63Eb/YVeQ46hL9hBaflUZaZqxvYi0vX+Vq
1XppNTSs7nkPecLQ0HlN+QZIRNayXVQukYWyvZsYS6SYKL/PVvK3PTLo7BnAWwK4SP7llM6mE+KK
rpKrXgRj5BE1s9ZQsEbOSvYxLspCLxQ1mczS6t/PIl9vgUwhh5LL0lJH9uLWmiEc1bF0c3y0cpkg
MUMQpsa7mBs8t7hpZtXHeW1LQYXC0nfbA6qU9F2f9AtaLFV279UMvPjzXDl1Z2Qglw2/lPRaLoAF
Mi4DCEjREUX/+8hAswWKxkVCog+uMFdVLp1n9FxCxzkBX1GJwrFf+lZnjyxQ/AfijjDavbSGxJKJ
WzErR4GBmjncZjOrGheJ+2oBgva2z4yZT5+NyaI6HR8KEZcD5XbsfkQy/QSGUCCaGCGCrF3goxLo
g4cefWcVQ16C7g0wXtwZkWnv70bJJ7DEea+gP7foxG+epSYXKIXpfYNLJzgHCr2p02FQVtvsuj3l
2U75iH9U7hy4O9IunIIhcFf8JdSUhL00KhTk5PAEeh60KMwR3IRnV9w9eb7119W47Z3FbewEPiIO
97kFeYdhRHlI2IjqyYZqpmy/6hpuAZ+vDRF9Yw0eQcybFKaFErOGTtfxjLkZez0LlHH4oWkh75CY
oCmbwP+k/UMupjVnCrmSqf9GM/WaRtCqWl/S4S4K3FTGSsuaMpbQfPM0LBuqvOOfUwWXXIQgZMDV
QLxxcAH6EDIG5GEg4BZE89h93arM1v5QlPYO5rPrbW1+QRdstt9Iv/h0Nz9XmTwQUgF2LkRzlKvX
bhUwHuwEgJOEiZBnA4eeW+/YAGwFIOw3H1kIkwoOB98djzM1dHXfykIW0DvQkw76D3Z2xfZt2riO
7PkMTqy9fUeMEyZ2Meg/9sukwzMdzCRhlvQGPwciYuY2/m7xUHUpO4+XDOKw+esdiK0pWPaXZTNf
BpstJY389fElCLVR0eU21d7SoIIm0paycPnp1IJORvbH3q4Cj+jrK1xr1IT+BwbXtpX7eDPlBCeq
U7x/0RK0CDxg+RIyyzcBQsnEHs5VjLCqvc9HIil+CuY6hre+eT6G81GVHkPxykSRegGERh3ZeTd8
mY33orb6LUxLzQvYRte1Fl57sXnYrEeKwYJgTm4j2TJjTXNwm0KJh5pULd31bhR4pyJg6p5cptk5
a3/F5y/b1nOuFcsjmJbVwLS4nphBOW3HxHWvQg2swG7MN+ilOXJ0YjSqr2HbXTJBwSFNR9fkhP3l
eboYXj+tb6BxXKF2G3gL7EwcqSIrqXQmV7yNW3kMW3FjjUwsYDWOjepryX2Iheq0UuVxX+Xd53Jq
CLwtA8TQ9tLCCSa4zRLJ4HFfSCpjFWNRtjzybqcRGQBz6QNdBOQVveqBlxrVNXR6VQzHim2eR5HT
sll2wqN5/ah5IFYKP7KbbWQNT7DztwjSFfCk7BJyRfCy3nU40T5ZvgCiwmkVOmCfzo2RNHt48sU1
WiwAftt4VJAlg+OCOHj34yp9CArUUUP7rOnrYzomi5U30yDetSzm6vG3ZQgV51Ggj3MYukreMVvO
Njn2kycls3VBN/S2I9a2dQQb+oFkQnEkPUP6u5e7jUpHaFxX553cnJ1zF3tWwkt+Q31OdHKWwEAq
GxASonb8w14v8dh+8BTDNPUxHB9zUKOUSkmp0cbN2tM6IQpBLXHCDIq3YEjMomtNLwB5u2ZzPWBG
7L+IFSdfu5HTeQwsMWgx4B8larU69G9BqMUVzaxpp9CSCfDHlFYcuIch3dxE6kF4hirGXfXK7Cru
+1k7aZPiOFsCSa8ktItM9bYVDetmnCZsRKPiEwp49v0/dDmBytMJ06DEjxJKvoOD2n9+7sENlh2Y
K/vax7Sb0uLwQg8PX320QCBClvi9ky/I5f91vdHLpazF1g+6NlrbmDwiOURy/BNh3B8TVblF7FFB
6KscW6Bmj8A43qAggUfK9BYizTU/vSj3OC339/sfTzYuq8FuN0BPrm1039ECm72ba7iQ7uHQyYJs
Fdy+G6peWGm3fK9PnbuGENZQb42XLifHnBGbdk2akbOG57bU66P0skk7HLEFROOffl/XBvLfAHMs
RvHaqs68fcwN9DQj4f4j+KFnBeR+skzxNon3hhzAF4r/gq8gCf/Pqdz1uPV9yX6fLV4mAPPIXoa1
/Sxg9xeoxVUgxYbsD3wiWtUJdm1uAU/IIeuGxOQ9nhVN7adIy6O2HOhDwUfaJ1gHD4EtjiPhkS3i
6p+lrSAt+wpxSZEIlAZOKhMC6hpHlvW4MsxBkNh6m/hjBFBQrR6AqaR+CbM9FCkWDWrOVezp2ca0
L+JnTTGdt8L4DY/yTpRPksUTxhLh4dT8n3NPsKSor4EBvBeHaHD+MlwtMd7d5wc9lvKskZ6NLSvd
MKqm7Ux5YMV0BrzC9M5K3Fq0U9I+7UjpbeePZgumIQh0NzW/XIijSkeXTeP/vg3QZja9/g2Xn8pN
JRw4aVwuxAWosKNfKDRVDH/lYtlbl0DyWs8fyxzoH/21v5Spf0uIbdEjUbZu0JSARDhOLZu/2tot
rsFM2eQDFpfJ5SPwyrVX5xhBze65NoTD6PXaOZwks4llbgSby6l1znpxZtn6ZcNBMON82PoP+Z7y
7B1zAuxtnkxU/dw/9yt+Y4oLYitS8tOXKpzKezpph3KD08G+5Vuoy0/kDztRZsmVpHrz03wVirHX
1l9n3yCsoAL/yBKaOsKV6ldOte6fqzdHoLzsAJ+sjHOqg+BMUyoGii1Pb2YX2bKY1/BWZjr7sdih
TqwzknBlfwl2CxqMWWwuI+ba8ZWWpo+iGZWUF2Rrq16pn/n5j5GQZFZsIwr/e6K3dEGW7Jpxqizu
imiqAWePHb5fqODoCxY/+IvJw+6T2bby3Z1yRwaazmp53Sd2G9ZqJxRTLF1p0M1AyHaOVagfHkMd
LRVPx91KCZQP77tFC0Ldl42DZVFLSJGgt+a0VW809NiN+vd6EpkDSrCsm0TrtiahG9MhIPHKLswG
yQYptNXslw6rYYVHd5ZghJhmLNoUmQAJIRLuESsynsEYM1KwrVjF7gVhoS56cEuxUdftRUz1EWl7
kM8vSV93BmS/oviD5ISZi2KHinqJvW2hw0IcfCO+lCJIredfmHQUB5hylUkZAcJzNcD22+z7fWLf
SQih5wkFvUCNzX8aqJUwll4QS3ns4rN1NRUtieQO+n+ZyFDqA0UHqSZLWy0Whnal/nSKfpxyfqGn
x2tLonlN3z42jRdRxzzzNhh0/ZxQ7AnSf1EqukFHjI1RSqoHSLYDKrrN4JPy3e8430otVGIA+L6s
FsfxbRjrASWTQVSeWkvC0sFwEprwNlZULxmePzGKUVwgXB4daE9KUv3+4AGQ9tXJbbha0wRrjpKh
E32QPj9lHJ9UyG0Bf+jjgYG1Q4uKaAEtBYXR5skwoTArsF0VPXc3R/7IClmwhnKNxvVdnxHpp4/g
ijIeBeQ6iILfgZjM32h+hA7VsVRMdNitFFtLMgfYeFWqiAKgwjc23pPiE76FXusQ822ufGQHupIY
LWQAW5VUdoJwtbbwC1V2qjCna0CMZUg9pg68C+PsGVwivdaVa+k6QuG3KKALXFdaQ/3R0mmY3z25
vqqqX148u8roUPaCsjPBu08ZbvHXXoLqFJmqobwGQdPMZ9Dhz8Iyn/cLriIWlpiTsDqCebzst9Ar
HIX2bqQvL00fz8QkuKPpgKsTWksWwoGur9lNMhyXUznJRmMrXI+LKOW068gRvLODgUrzQZwEVety
1Y6U7UWvzWbRNFrlWdMrMlVBNXeN4uQao2Q1rldbXtRrStbfMOwYneH8FX4jnx3h1o2rNnTtUfUw
rClFKTA5jKc9u72w5B5/yRd5flMA2cljovYikx3pEzf29hP4D0FMkPTZ+7Zzn0QT/nqQE3/zxWFt
TLOLowRQvwWnKCCcXBHaQ8VLHk5daMRCuD2OQnag3NMo6FY7WGhjHbgKxqXVg7EjJK091dfA8NqB
S6Ry9Ig5mmLknISxlaWS/ZvxJCTu/nzKPIxhIsq+AxGWp6BTD1VBG93qFkfvU6uC/c2IXyT3nt/d
xHDWQH1nDVUw6hdu0gESqGnPU0i14AYPUhiZhgUaB4GVOiyJR4aEDu6/n0jj1fKJbM5lyiRqwJIU
Fyzf9dvEsIZwMDaNXgMPeNneKGR8vve6FE/D260Qs2b82X3RP15Bb37EXtkujPBSvyAnb23HjE5I
RKEU3geCNQxXWZMjyrXXtYd9Ek1j0cSiF9QkCRK6I558FFzsCTjsY66sijVjI7kbfLVnj4AnJv70
29SYjA4cBgyQt3YttB7YwYZk8EdGZNEHXYrpLWT+yjmL/LgEjOkqn0OMPepLcixvye5/u33sIoPg
SFN/hxs57WhX8oixiJNlOsUCrZWP7vyjhJCAGIHVvuDK/6CMmBZezS2SW6/zL62DjK7sqasIf2pV
Oqnn+7rfdo/HKalDZ1T8lxLJUOlBl01tzF9igQ/vm83DG+fj7/7u6ny4X3PuLBzNYi0SGejG0Yeg
r+FrCeuAi44vmiPdUOqApuhhVy0n1eOoJ9JD+WZB6Dyd+RS95+mwugoEuQQLIvAD+Ub6UGsROmoU
5U2+mzpeJXQg3wOvwY6heD7TsyHkPVTjzUJMY8BbWJCa+jISAY/2PIoZRqSOQtzVZtP0orKolV8F
4Sn3saQWsr1rogiWhgjfUuvTCNcrEVxWDDjHkugu8v8u0+xbvdkvRdS9UIOuwz/AmzExJRIthrmC
cm106T9eYSzY3AK3NR/eeYL3qpOOxGwnFFDr0V1p1l+GlfT8PG1mSBxKry726kOHKOa3xQ8I6Snb
cRwt5DEPlmBcBlKCe67alZX2cYMWsiUFdjyo4LguArA79M+v75X47AOnJ/Aw7RKJeNo1b9BDZ1Eb
jpJLwXBYmRdSbUBRCyYBdK8nuLb736eyixEfPk2usUv3W0Tt1tYDnsNdvsUalTzaI92A4QZZ3oLy
vy15MPZEjc/EpoaJYrj61SNn1FWat3cQ4ubKYNGg6BlkYfvQhMu7DeMIrOLlCpgUwYXUVX+s+boz
9RkDKygdGxaCZcq02JgDoKdj82TXsbFMy5uFfXqe3aC7Vom6IfgUI6s2jHprYFmI+RRATr3xwWHQ
JYZp79bfnoMVf4AtjCGUP11HA1t09CJUSTI3XCxw9/or1cs+t7zsBdEFvEePhgMTLHlrDuaM79J3
XRVI7EwVk/2jOdWjcgBxvvo5IgZVqKIxQmYhG4hSuIgdaF7t/nXn0Fg9t0bkbQxL7YPuv19zjMoj
rQF7zRJy+BM2JzBj3+PamcKPKaOHFGVpVrULUOfXg72wPxRJTJRvEIryYUuvS0j36GNJB5W98tlL
ro+z0OsNWND1bSWZUBNKdh6aU+q9pD8ym+eh8Rh9JLAVkGjiO/VEel2B9cx4/vRcqoJFE6DNQv2j
BHsGHza8MU7QGIQWwS5MRI8fwadTXSdOfxPpDvQJoUbGDiQ7+3y1uf4fMcUye39NN9bvpqMAjD+V
+tmZXLqr6tCSKgkMDUWtv1jFC2/rcsP1SXklZ64ze5LcS6Tlh4pWM+GbcQewwldNbUplzoJLVowy
Zl3tO5pfG+wvjy7xPzC6LhyFTkjk06MPiy2uT3b8gKhN2h74/pjMvMWGGJ9Lw+USYHcqWtVQgX5j
4LQdhb9OsVLR2d3YomoVCz1jQewEC7tFWNZ+4IusYuM08IsP9nO/xPPYqOh8MseoI4GAuCHEr4TA
n3Utqg2YhICr1oIOS1nrWBvHb3aJMLmC4SEL7g71nziQtl2Eqs2atlLMeNfCLKbs/YcleZkbrarC
4GCVls+Dm5HxbPKbqfjiVQo1GT0Nweiv1srqDLwSsw7labRCXWbmjlANOGw6HPXk5xFl6Q/u3D6n
SbJP3B1E9qbby2MMvha6xqXrMqkXVSw1Qr93VHJpylCC2erYGHMEPd8HYo6n+G8Bn7rxH20EO0Zi
jO164XAw2dldbLJuHbEs9Ap72DeCWkhg/gQ6mclbSXhskEroj8Pad31qYKCkl54qgs0m5GAwdH2q
fth53+0ppgAAmPr++IFlUQPFwz0+ddO5MuFQbGnTblnkPH+1HQiFv4OPm2MSMbjtomld5HvURAF3
bIO9SXqphKc1qwM6Hbvg9r41WsZgARf+qN+F2jewDsrhRhcZiKOvYpM7EeilW5Wo7XJKIuxmATjR
nRpceW5vOz9dTbVXMoRxuJYMjURpWRi/I6rRKkAZeGCym9b8h6iEGhaN+ln8gLeKrbh/SCSaQVck
l1W/8fzN+GdQ+u8Vn8q+Mll3kIxyy1ZmMSJDDzRAF008PNUOttSJZ8a76mbluI1Emf1BcjECKbNn
nMcnFsUyHc/bGHW6HrR4xRAo7wootYWK4XymZcoKU3pZOKE7oV5sGjUMaWKlfRpUlqIfvl+ffV0E
jtazJ2i8b4YQDIGGMPWQCSeoIuLthXuYOmJBBM4k8DXpI+z9LRPh5QsioMQ0Hw+rwpKctw5Rnf3z
ocpkTRQnEgIxyIsJ9r3pjRYINSLqr4TaRhmT1rkmS6zns8ka+ZBBa/cHaSRpl6O3htquuGJkJNWK
5EJigLRtzEgFT+zZWX1TOh+1uIXzD7yh6sgMxNmFXhYvlUBVN7sZg+7X3wD0nd2jtFjHSQka8+RD
/Grw8uVVKTmvc6W0eKtVB3qPNDsENckuhPnvV5JwVnLtNGochISsUjVzjjGDw7k5qwFdZ7ph5CDx
i+sNFuNbMvILaqmNWrS1zMWxwcYxFtQKkhmbBjen2es/H+wBjLLO1xEqJq69N2iHNnuHfHZVfG7k
zum8WkOX0sIrgctVbldNrA+7oLaYl6TldB3FdBU4gjdgJMmvy3U35g+4mVm1Aj8Wnjp1JP00eJpb
1PscWf4x290/Vd2xMljvT8z8mxzL8+ExVOYsnqWOrmIdgD8wuwkC4xQQEIqaGkCHw/tvjTfAhzAb
BFS/mziIjlIFYpBz9rc8N1ICA4NM+cQBAh280CrG1/RS80PJFJB07Yq7sehDhiS6A2muBYBEbODu
+wjlIR1f1ai0gLLBeJkk8KwP2+Bx1cdZU6U8NQnbqsD/sQGBpczzbVflVlhrnkmCqxEIxWqiMI/1
rzZ1VRO+zABKCUp5C4+lkVWr9k56gFBdqQbmDGtu34jq5ZH2ssO618lG+bZ4ozcxA180qtfmSRXF
FM7MYVUwKt6WyhT0kf+EFY70RmlBgCRCbrkAuT+IP91mdLJskXWsVpJIsMGGygzsxxBnwYKeSEVg
q9nW1OZAJPBprNc/w35JQodF3bMiVSurx4rBIK2uJmCivEkUaYlkiO3MUcEtqaV+d/6DVFEZbzZ6
ZS6qY8rDYhVu3dwXcif1+Ao5wd1KKbzoYzRrWjN6dsFyMXGLXl90kh6ke+sUQJPO+Fm98m0fm4Xo
l6+f/2GIHWr84nsRPkXmC8Ljoi1gRXsIfT2jUBjq6w7n/OFs9Qk4kB7/CPV7RNIH+27x+l8Zuwfr
hcIZr6cXZtp+ozYi/XdYDlFOpMiPQyQ+ZAL6jSCTi4pMqxB1+wcL4ZixyFmHyUtT9AC73X0A+fNG
EizUoGukD0nbX7XstaUtZclqlhyTtXWMCm8n8A1wY2sJbC2QpOYUjesOF86a8pKoMI7Xf3NmKhhR
/+EmE9qY7aPlPk6QZDCEwtUdc8PfWPwQdeYK6GMJJ2u/TlVt2ft/OLwu4euWTZ5zOdNlitZRpNbE
1YdCoWd/E87CDS3CcW10BFWtUl6Jsvqn+iYl8rQqVtS/sVNwV6A7/1NEne8eaza/6yEDj8iOWV1h
VcuqrnC2lPzHMH/kNmiP2P8WXnBaomnhiv74ycbtGL5eSKWwDI0JqUQ70ykiER+Vj7l1J0Ao4R9n
lxpf4jVZtcVDMACKcgWgaR5BhWgcw2ZlWDmD/2JsQPr+/A4lAye4RLIzpNImkYoILK5tC5qp6/9I
RivLV0ycOGo2btr6Gs1I0hSfcNiygAt8sGBuK7isY+XUycfJt7uPfEhAcYQCpxRk9xBK4pOTnKXg
BrGZmW1jxNLzo8bCwGXHkEWBecyRTmwB7fcjv6GYDJvyKFhhj9GV8L+7alt1inBNjBbQm98mG4en
wAWW43145fW87Lg2lgtZUIKqPwCaIfDxIeUswV+XZ430tkX929F0XFq1q+2mrAsjOIrSqubjINlz
mHfJHqijZZ1IhbpbENvOxTORXdF0vPj/zXQuXU20ZL3EcdVWc9+T14jK7vVX9ueEER4qPkFlkl2Q
0mpVfu01JynIf3NCq0kLCS/AImR2gaznPagXDM3E1xSy6L2108vxi1XV5JbgMaeYEs1YHd/FffzR
6f02381Ccln80sRh1+dg4uMczWZbPNQ889a/g/ClHIa+VR1BbM25kr0Hd0m3GJW67IebKhlZHY2u
1JPU92PBg1Plxo1DUO+4hnnCQtXycH/eTTw45Dg2tbDxNPL8hTKz9omsA4LAKyIq0ZeAkXI0Cps6
5ZDDbKTUfiv/UKhUXNDQWs8nUwn8dOjuVCxRadDaUBWslP85U6Fgxu+RymaWL6HEm2P2vnR9y9+h
rwWfHaB6/DOANWe8YG1s1K/3Z9c9Dfuzq8bFipH57c8ZLic6adM2GFw87QqtBRTRTFwQRLE8gdV5
Jn979EYkNI0qixpTYTR9sWAw5OAO6UwiAUGdUnraQkJllOmaq3iNcOT4XGnSJD72eqO0Dq7DXDll
6szy2Ml2B/jGdqkYiTJMS/FPvVpuYuitfx7h76AZ9KPWe5L0X4BxOAFd+Xhi4ci/M6IWeKx83VBv
sVBNrTxbXvvQv2cvcZ1ze3Yjj1TcwPY1QW/7/mvwpd3GMNapkP8zAFOS7jUBmH1O2XvFhrzBIqgp
BAHbVhLrw7aI4vYKqVFEqvz6r4EMhKb8KF3ubu0nKSP9UwGJ/N3IMwdLlbAhfQuYcFs0CrXn/xUs
QXUEI8/PwOm/V9+9EUR798ojFz21C7aLggLXuoCC3FvtuKStf9JHkTgaH7WLqeef/DGNZ5U8vlGv
7wzi7FGkRBfz/nGIPFuECfgyTklQaZloHYLrHr4DVmyufxIueWzJQ4J0gdCShoa4f098EYV6w3L8
O1e3wTZcc0OBxp7mH1JgfwjEhNsM1/J9S+j8QpSVIipLKWIQr/f8AXkT+19zAcU0uxK+KQiZmxoK
wkH8WjkOBma1z84IKvJ80Ak88Vo2f+io10JqVaw2qX7jAMz1WB9Mu+Cd6hkkMAqgUGWqfKwy4kVb
ZxQpixLyu/iKgq36cEEJwvqe2CYWSpHW6PRFqI5ZE6I1fZEYvgproUyqk0W5Uk1+KiLLx8prmDDp
oVimaUsgGOtJ3hx6gi3ObucihkoDEKf35EoAUy3OvnfSv6QI0EugcEQ+d8TPu9aYnNZzDpohlBm2
gwwUFG/zStxP+w0Xh2sYtzfPUPyk+sHHZCtGXUD1n7HVrMdbRXs/zAgDSwnoxaUyg9OisPMU3L9f
zPCLRFrnUI4BYzdhIjJJJjicSechQ99gJwgwyRSGN9sFjV2bTy1HIoxHJ2rJkhHKJF5Qua0tRqSJ
iDnq05xMChVRGEjfvk1F9oss0jh7rYDmT2oxiDYarVyRNUcVLYU4M4/ezejpXu94JDQEVPYbvQR8
9pyRlKagvp7XlZQFUwIXJhUDhKMLSAO01Ilj8X+jslEQYIpsnqN6MWxnxVHWpaB6Cy7IorsASlSp
Ncz/5u3EiLOi6zag0q5kGld3kz06zYnOW2VpTuCHgSe0/VExwOBd2diWTHPTtAzx8E5hblUu5YlU
DyvIkXwICBsU2PvFOOMUT5ImGuOnoyTBv5lvxpGUiHbA/bO9/n1/L3/Xst/FUgJaPkxEAZAnXCxU
x5y9+7lqxc3C2e0iyDJVzubt4fQTCAvMzKq3SraNYe0Z9ECICwo6NY8jCwYTBIqCDqkal5WCteNr
U9JxxJVUR8Mwy1EOA7uQDtzwk3is8R0w3Nyqz6pMB0ZAMBL+e5eSvkutWlvHrY31C0SkOhslK+fR
qHe6a9+oPLTUuDEu0C15HWu4HrlKbCbvn4HdCJKQcr+wJE+JSqWNrjJaDwnJM6KFHgRxOlwWtFM1
gKRaWMGwcmCFzh1IrFYMcD6QTpCKamyQOCs1kK81yBgydTmNNVmUxFLFlHuVJ2mDcQ0NWBqGbF5s
6ybkyZBGJQUENEMAgiOINqvF71UuMnALKNh+8deQphQD/g06bxojHw0jkywoHq8vL34E8dSdz7xs
Rt2Dz8Ob7rnS/5zAs870oLMrtM6KdOMPnBBLCgRD7U1j6yUUF6UxOEd0OiNRtcYDPpd4vzkzuB3D
ivGaNQbNQN7bzXxiFRoiMgpH3VorXrzddBZBJLLbK59Vpr71qDtNXgZ8nZKhW+nQxPeEwK4u9WzB
XNOuJbJvE0dqlWpNV1NDCQbE04Q5wgnDn6jO6Dfu0qa0soOm5B+E7TirYvcU1DY4YXQB7uSEC/NP
NIzQ4Znykj0xluMYZ2E1t7nrddLf8gdQGPrT2wcGI+vwV08GJvMPp97dxmwmVgbOvbQa49vZYTPk
di1I5o3e12QqCUclGVPz9YTuiAzJhcMfbnJRa4vdhrmDX8pCaDsD3uJV7HU5ldPfZzXM97tE2zqM
Dwe+vbKx4HVf2gJVq1MOd2JUxd/UmCtHoQgb9oE6tRWj5DzDbZke+XJaeCIbMuEWfN46uCVeqmu3
fo/vn2RuS1uZe6SvZZb27ifyn2YfXpApXCvbDQATvEokrJsuDXLrFpYMT3nFTq9g+H/4eCoGqRjp
LwBwk5feb+Dknoyh+hjeqCuv9g/M8FkdnBP8nw3cPnURK4s9nuE64e0t2qOr9FcKZ2xvZMOQrWHM
kSOU8dP4rOC1GB5p6ObqKibkY32HPn/CnG4ZXeD8YlcVT2WoYI006XkudSm0AdIQHL0giWjNLre/
/fjp57ovfuElzJxqhXqiizc+fSMlOhqnZ4Cmay2P2GRVIHrF7vl5tUFJNcxieRXtMwpK1eYkSzri
zSYRPPkr06xtYckBuJFuqYcG7lptiItSb85mBlTVJcLSFGt/gakLBnnV4Fzk2mWOpx9+hHhOwSmt
ZFlJyoAHjiw0ySrtuCU4IMckdBPW3xWsD3wd2VRMdpPXFJ2AwILoThDT5cj1lNJ/akxujt24Ys0L
wYGqkIfJLIPhTELyPStgv4NcgNREiZ5cue3ccVpuB1bjowRUYim6zdkUdHIb2dPWD4NyKxU4Vrh9
DY2L3Ok/7MRjn90twkQY0nP36IBGFjeErKUcORj/JHcg4NHT3z3DuXvSZdZIKut9msvrKg7MWLUa
tPl3QnDLaYu6MsW2IKnYchuO4kwT8zliFdMp6PM1jTFCggPgnyzgZD6no7Y9/nmqHpD54K5LGLY6
1Zbijg+mEQHLwo9tR7/RhYNkx44R532sEAmutdse3AmTK8/73cMZiYwM5vDiTBIlYvc9rLSEoOGJ
VLvWdi9ccnqZSRnD+yYrqWPtwQ2F2DyYc2SXrHUfieRLe3b/lYY1GDw0twU68L5jfM2DEUsWGdl9
wwV882zwO0Eq2zmhgErB3UtbNvO0O9Mp4USmJhStfw1mj+bfs19Ot85TpK+o3pd155L3AvZcO4mW
yN65iUfZwBZZl8gHhc/IjK1e2mz4jRajr9fUFa/gFPwO+QSKYjnaXp8vkDJrT08CK6w5LQL+niMf
w8usdx/f7rWtFvIXwth3FrMAj3bYnWHLXTFbQU+qAGl+MVbHgm0z/C7sRTSSkAiHtXwyafQxOGib
N8qyIBNwXYXQppbnjgJIXgaDobHgyCHrGAH5E8TiDDfk0SOE80FF/i/AmKaPwX+haFDJ8cQC2kJi
ZNsMNqCAy3VMhDegzLzXL2FL4fx79YC88993A9rYZ41xMv6faTOXY0qnG6d+nU00TnT11aPLy3yk
XbAXfI7S4Uvz4O7zQeuoWlVr6yOkX0Eiw6u1iaNx+4ybOrqD0WNMCE7iePCBni6h8RCWkPJAvUNK
sdtiqpiBGfUSF/lYLerRdP5Jh6z7CmzAlg9GRd6J5q8D46E1GwIteKcdoFTTz1sAYdfHwb7nU/AN
zW3Ge6vcuL3mMn0OXe2sWHK8L8qFxFJqqHAdqhLMj3fAsz+Fam4bonxL7qb0rW/HvlSEAfhU36E1
QgqHMguhhKbWgbpH1F4lrAtlY3oiapTfS6yBq4/m0xLxFjsstuuSxkloyVpGvfd8zbBTiba0ZyAT
UQBCwsZxXIjliaSPkfTkEmqsP48yYi0FRVRCe8eg2hAW1h86gKN9tuoIq45lnk6brEaRbkaOE/bg
lq8ITwUfIMUki7o5FSHZuUgCr+qqEn4VZuOZjn2cULhDeTTc7uzSD/KyqHrCTgpKMcqhiMyCVVxM
RiCHQZH2UrXtNH233XvLQ1yimji7+IhiWnsVLY/i8G0RXHAYkNlXm0tGOJtqfK/3md4O61eM++8l
R7U1dToOLtnf7rX8Tqbg1+O7iooy7k3M/COqd1rxvbrFzAaJd6cRVgcXTfUkom32qM+wWDlyBN6s
l9Qtsz/xkefRn+jEaA7cAHpggGGEE/wqVfRfA12jHebZOiDECgKxRshGmPllsodjl6+fO+ErgNx7
yLqXFs1tkXwvXEdl1RQuuCtib98a6WvdCIHi7DhrYkp8qIhCHQ/sMOP2qwDgTEP+omCXUH5ebQlq
U5nzeWkLC370cjtv9onnEHdKJZh1Pa9DAAeIKTfhb75X1xPJKZEJ2SabsK/duPXrrQ71wuSJWW3d
ptIgWb1oLZ6rb14iPGMRcRGa+K7sEyyDwuKMgZTyc52iRzFcTFAzto1y8QF39SgwUCiDbOTD1yNd
Jn/2u0g+WHcVsxd7RY9uxexB3qnX8eKAkaFBDVORyNALhzfy4vDYIvJkcxX5bQCh8CHR1rXvbp8i
9XvQSD8z4lN90ZuU5KouvTVfgYgEpYEUAHSAqQ3+n/6/QDt3P2kuxF9zGf70/gyHSq0ZAfKF1bXV
ihjnFB6R6HhPu/E18zwi2jsU8IDfjeann8hgnxmSk0qo/r5JvBwBytSkPPB8Lvv5QgC14DRzANvr
KsR2ADE6gaK6YmcWhKlMzaRR9hSvyNnInCIIzNcA7ihKoUMlJg/O5dot1qrunQRHtn6X7GLn1Ijs
j2Mk8T0+9/7/tjbUvkvlp5gel9IGYeqBTw1aKt5IQ1P0mNqsq33aercFxTxlVmKO8wPm0KhfgVDj
RFLv4xj7/nOJ07V8AduxwuQvARDMk8aHt0eLWINKBJK1VpSFkD1yldqiLG/3oooXK4agPjG7qIUg
IjnMtSGZI+BidIVI7QsmgD7dLyGyMEF3mX/faYQRlzCtavcX6LwnLzYysZMRTqPooSU13MfGo0TC
fTWaWQ/kyXxUCndTojbKZZMPOIrHN/WA0fKoJtwntOHt4iVHGeAL/6ro8ZG+LWNNCCFhmvlsoDdF
U0RIM3atIBqhM9dgUNXsViyEpavpipxUHHuwtzJMepPdPlm9cCqJC7kFfyVeHuHdZKeHZzkGx1PG
NOft7zKAfAHTdX+WL7yL2omOPQ/1hLNelZx3kHK9hD5AqYMsrOQt4qAj1vBoXlY7YmC1BUVxjkBq
73rPRrRg6ezum1cCMmufSK7oh5qxz7y0sGrrGvYgooxmIT8Ixmua6YsyR0CkiDQnSb+W4ePUWFsx
1tvgKBTppmLPscILEgKpaeE2Xn+uubz6bfTdvHMnsxs6mdRsh5lUEsoW2npIbUbQ0DSWvxHp6U2Y
9f58XGX2omsby9kpOi48P1ACt6ojTbECYj3DNz8lp/R/lxUEsOijsVPzLLHIR76ac0ClmemP5ysi
7l275ocT5Wyn4PCCDH1QuprGyTa1cp5WtIw9VgLVsnW80oid4SELjbj1s6oCiD/U2Epu2qYcCFCY
Avv16JUZoE+H6bb0dym9E/3+fHOSc0urHqfr+1+ppj5QpeCAT2zwKoeB8ClM508mrG+mlXoI7oAb
jpDJZ3PTH3xtHVvyo+G/DOSkNfdTHdXVJj5fb0X8IHnNtW2mx2AeJvfvQqJJ64bzxeDD050cEOwu
RCAyrvRJhoyP7WQkJ2DwkkQC7BjC7LGJsLj0dak0OLh8dUpOoF3BuENgonLfVmDd9uI3FAFF0K+o
exvx7CyrtAVS3rb7sTIcuXFsGVvAz1jCxq9+0BbElpwviU08FfJyvr1aAzP4grBJAU4HdKTlXDNX
6xE5PJdMSly1w4bcwC24ja4ieQ3FPFGXp36Piqh644yZCIadiYIi4FxIKiiE6eIdu92AUpztbmz1
Y0GZtHHvG+zAlwUNOS9vhMLeun/UUTzY3CCW7uqISIY11tSUOKzAfkhG0PqXHgD128oEfm2JIyNG
O0zq8LecPzCKtqa6daiapzvnIupqxPxcMYbYZ8rWVpZyMuj1t4cC91U7i5XqfshuJDBcP4dFmnjV
pFHwqPF6p69+BPTDIxDAFsfhfyJS01uh8FXVrLrMtbmAPAj2VMMA6NO1F7tjYQiv40Id5NiN9+Vb
F7DFVp+x5TVyC7g4OGsIwgTQ8pIn7GvpzRt6JoUK9lRibJ0DPFxT5XnuXE1VYSgX3JdvJYRz3tHR
Z+zXz5j+2an3pqbuh5ILvYECZhxAVkVURxcdWKI8nnI1y8ZN3PkZhwDiouHY7je7GpNa5D6Me6fV
UQ2DdWZidt3UasXJKO00bLbKcP2gcUeiO+z/VhPL1aZkoA0RRM6ZPShiRbO5+SjQyH7AqNPhFPUV
7IJQNbDxXCqAew63KcyCpZmfRPo42Xww/kWgjlnhBp/EKGlmaZdVw9/SZEDCi7sW8qs3/zCETBxT
1p5ijd2g6p90oK4g9MSxZJ2VLBKOciG3/3X/1vpBryJozFh45z/jFOyYhBmIe44ve0g0FK/YF775
rcVdWD6cHJD38GmOVM9v2ASRhJ77P/PskQXizw+BaTzNg0NMJ9VnfVjyGEm8sR0TubCnrZrveQOa
uJffUOizTItSLUMN9VFndymGPOb8mASrSkOwtj3zoj0KbyPdgxjRBtB8+6bRz2fhn24HSjooOChq
XwzE98Io4O+aCPRVjHqM0C/TFxzoUkSteS3SuJ6DjE3ugx3t6yWArhx43CEeaVXu+jdnujeJ89Rm
4c8lLX+Kn5q7dCcJbsL1S8UF36t0ZUzzvELOjPjnp16cVQeSZrcmHIXySJR9ymBzLL17O5POmbCJ
vIzdC/Fa6oZj7VuaUZMmDD7+MbKyHqrDcwhMRa3zC4mGmqwQNabVzi5LWddFm3EsiyG5Fe4gdllr
IxEIysJtd2cKRDkglmwuABN/78KuqpDNseJCrsZKxnLuZxhY/Iq6vtpsKBGUFWptx/YxEBCxngBd
vWUFZiX+UNRmKZVxWkcxmJHxuY0SPSL3E5FCfetYJX2Ia5NOB9B9TdLy5OPiVSVJGbp4CB27WkDn
/KA2ma+rT0PPn9JGbFLqK7yXOIHGNXb8k172aI/8/31WTIAjHpUWAGyIcAqE1dbPYotLodY8GrSh
J2PL6Wj1/cgej1up2eOB47Qbfb675lGSiRwftrBvftCk4Zj86lMm/SpKpBURMQdYZc3Gi9KpCdjG
P0+QL1CakVz1GnLZg4CK1z2iJr0G6mTo+XGC1loeCedIbilXHkayLncXlumnT5f4jI4MUVSE1pRF
rVTQdPr1vqNGzh/uzp0cpj+P2RvE6gxJKeYW64xf5zV2t/p6O46bezwDk3LbQKRyMWYLKuWlEt13
GgTdc7GsrpA1HofEd44AO9/RTE91VnULoLAxkkdNB+5bOcymmyQ6QEs7mH+sBUuSEyVQFoQlg9sK
16KC6qu7uTlShludLDa0daBRNmNas6sn/ZhdQnfbGmEikwnUkGu0D7fT+GyWpwOGaFxyAx71FRnE
cHgsgN0EgWQAY+ZUoSltwKfC+Oz+qkkK0QD8u/ZNCBkyzpWJjuy2vrVFgyNF+aketFlT1EgGO1Rg
gbFMmm1HGJIPn0o+Qk1WrU/qmossF6gcLwfY61agqMv13no8AdF4gcyzpMGlr6bRFEJGMoUOmClp
zFzWs56E1f53fOJ3HT/3J8A0hDOkW02bdvt5QgGl9XCPBiRkHhTp2hNXKmURW4jDgagc+1kYOqMp
yn7Q6Y+R23Lrwg55lznQTnj9L/8nZfmS+3KsFaDlDn76NNywCKXaCt9Xp2kf6UAcCHZjwkhWdIgI
tNnrvqA3PDnXsJWbyKtOudag456S0Tll23A4SiV3iPuvfVjWjeO832ifStLhAyEd8O8ar2OSIoie
e3bb0pPoMxY521qIv3mWRUBTZ4tEvE5nxjKCjx9CcPHD4eCeWVHhB5kpAYlBO3xDJGKCp5ZzRVDI
t2RbW2s75El/c9oRMVL2sX7lkmUp9crFDFSX2o5DDWtucenI03ZdcGEd8O+p4tlbc1gdtTxXdBRa
nGaIzt/zKXLBAq+iCyR/rF0w3IV9yY5/1jnllMZu1aDaR80U43q2HV2qmKBJJsyImL8DAvdcXxnA
EZm9R7WisySQ51A0ThvX23WeT3MWFulBDNcQQch4GGqvDSp8ytDM0AtYTkIaHubqSuN0/Hrli8SF
1GesjoxOUTNs144OdSQlBK36YbPXH7sHLU0GufWxRHJKp0dWKBDXv2HG5ebLnlXUiXaSTE5dxB+0
rGWj8T2HH4vRWNxcvIzdrai+IPzXMd1wn1S8RRi9jJlbIhKTZ/mDSw7JamcjgiqS6MKm1aPlC6D6
kJkWyvkyGCv9Uwt8zHwUrMLOaz8CC3UuRCXgNyD1PopXY+L9Re9ipnwhQZpJFzon4fX3JEKodZ4N
bKaBDR3mxvnCpCllcoQ6tQe6SJdzTkNb3Pa/3FzMLjNOsPrJf9PjK7m7R0N4/TT4XgGLGOVhonX9
5zC31oUI44KmaORrRW3CIUkJNZ+5xngq/DwR/kVIWDzoNYAsKjg0U3/2rJUfyus9Ywc7L0VIcbEV
zzcl1BWZstvGgF9YtEeS6aLYjauBKacmHv0mZoG0RXKEPRbxMdIb+MzpxTSW693Vfn4xECzTWalC
b3H48whj5zz8+8ahqbAiNvehrZuRDyXHECjeLm4jmCsaHuw4Jfbz6KtaayALcXdK1lpUlweBabN8
HnffceKWHkgV51Bv93ef3F+MfQCUm9T+P0tvU+v5mIrRzTfeeYnRJXPpicGXN4YUVemsIAr5BzUl
/acsd5VoOkhe1Czvi4+JVSc7P3l2KJLywflMWxxvTNfogWNAezecWYvmwI6tBORXJKr5A+bsVx7X
7vJZVxMmnyuKXhjlJ7GyxgW2z+rm3oLe0RCkZ+mSH9HJmOpVGaIwPCBOMyJ9a/cek4c/aozoj48u
Fs5a2qF1I2jIq7e+b27ly6FOiEQGeVScHvOgJIDgu7xC4zvS8mBOLJeK8tGTO1yQ3+REyZ4bCAsf
2O/P0kH3uBtwCKYaG1MfGFCYVAH5JZbXsBq0WqzJexYpfLyRo4IaRn+u1VbQzE0X0NTPVl49Raek
vhnO0rMChNajETlL2uvH/G6o1iLhrGdbuWq8WmslZjlSpCrtv97z3swwaMHl3QVsxf7VP0rtZ+jL
1B0NZfQ2fiAwJ1AoyWRIm1AqYBsVUQ8mbMl/bynx+pE2hQ5J/709llGvm/U6lFww6niDip944pem
le05ooN21YFvzLBaa5XQwMWYbBGTBNNZlTaxGDe4HcyBzWD7XwoXhBQMeintEiVo5FfbQ66gIioU
lmu+rgLrKVEKHexnq0EePJS05TcBDKBEqheMsIrem3T9e/6rGYwWmNnKfRXhTaCDRQ3qyqEqVcpe
WxzPw3FeLPNUGPOJLSEm1aVaTHpYbNOOKeQLc8Er+d0QaAW9osF0tnGKfbcH+VTXBKsZK+0JhRhi
xK1P4VKEYBNUsv+B9Wt1qs/omIJgyA3KxdgmuILNSQ5blni6YTVr0gtbeBBFPjre4qqEftIjxnJh
k82Kt/ESHAwUtXVKP32mA2XNELd5VDQzK/swEuSU7V97/bHpcQQCBRTc5bXgkquew8fd9Y5umm/G
59BBgKgRinl+C+Dcs6Uk34Xnw5uoZEAhlLIHzAyXnAlPLzV5tnE0ABQUUoBcKpWll5+XxYzRYgoG
TJu1yrENLdFvWYD5s3M9SvXcRqI4vbubKTcSVsuEzWdMM7ADMHQwlub6QI6ycI2PHPSXMoxVKw5N
dk0NMyq/d/1xBcy7YCNmZfd4VxJjVGdYHPQi+1l+xVQb373VdietrhgX2QhZ7tH/DFeOAPe3wooU
ikb5qFvPcdGvrIbkZgrEyUHMC4jBP37RGofW7U/EWCo/hlKeI8TIwPq5kg0Gz6P6OEBzu9WUlmbH
CU19Wq2zbCzcBtv79tFbZGqdOkoBc2h6FqXt6iTLc0+dsufg601sQea9zj9IGvs5cQklqdK/u9ue
KTj0ORJKoK7GYrv+ImNUSdQgm02p3gzsjyOpKxpjF46utncw5GlOIunghNnyJQX4Ua/wtDB8v+TL
LX5ee6WEaGBCsWplHaLmmpNN8fzn+VK38lOzsjNdiDloW8xzaFaoUffZBs+k0J8mUaFuxBpSwcMF
HzrLVzMTvXiQ/VmI9C96NkkUMYau+Y4kljs9XW5s+RPcnhmhrgqRRe0aw7GBsrwn9YVtYYcRBb8t
sFw7TgnzNh+ynwrlgpEeDrFycs6HhcEMnSqN/95L6WNnIb7SAc259Juu8K38tBE3ySZ1KkUJ1X+k
CaKQ53UZ43SD4/g1LvRpd/YT3GBdeXYvlIHqz3AonQVvCxngCANtAh1vv3iggPBeXqS2F1d5/AEb
5w8Lhe6SCRYI7KS04I3LvbaqmQyci694ayjMPzgGYn+6BZtmM21L/qiuFEMMRCjfz4e4zZV15ev+
f/eF3MWnBtbG0TuJMGBYBjj1hAkCDP0Qv6Ddo3lgxotBm+Gm349YUq7BWdxr3kGN0fJCLWFFfZK1
/vVM+1YwnMNz1SJ7nL0SphhEbVxt+kk3VFFuBcXRHNKXzq5GpMn/47lbBTz0ofEs4pK8S9Jmou8B
MEwEHj3XN5v7N5U5y2jO8tQX2r2Cl8u5FeRxtt4ADF01Vo5heG+eN3wDluY3PPFYAZxQX7Zh6A4+
+Wla0fOMTO3KnbsXmW1zhu5fVlh58CzIOicjkyKwnFTaGPNmAZD8e/qq+PRJmZbCB3vuHp+7FUny
ae/PjCAH/V40zNbbhDnAq7rEvhnl8YRTbnsX7VZu3lWKhwS6czfJKYngQtpxieZIRgqDHNBTwIE9
Jlbhrq6VZSAzRjXj0PQFK6wZ1fALiFHPhmI+4ehNG7r9p2hlQfHgLmjtzWIIZ8z8HtNuB4SYVTUg
5RgerZJnvCBwwul2kpzExX+p2o2XYKveGYa9tawW5WBNqJrMeVkJ/rkZePjENSNtdiH0TmrW+KIx
uemTdTwbBudzw60i2z1sJnV4xBV4t1k3e2K1wMcWYDD092sdXBifj47vIEKwTSIHR6FM5VAgW/Is
tcJlHOE7ae2Kf0MLu7N+7WalG6zeMmgbZnfkOc3I4y4jWVIc4Lm4ke1b1VlvMZIDk+XTurhjxvhJ
hOWSD78tInb5o6vMtmZSFVMkcgNtZiX7Q/hGmVxEHDaoe5RSZHyp0lQLGFibwVZb3dlGvE7GjH3/
hs1o+f0fVW/dgi9YDVHOVvJ+b4RBuv6620l881AgSslwVsgcvXj23J0EZmq+kgnOAs1JBDYMyXsx
vHUCW9AsUpSRlEe/IRs5R5lbvLrNRxtxx+Tc29ilngosmTGNbFMrQH8RhiFemzXk6NmFGncLqYTg
Q4RMLgCJ4KqD3rieOkWBgkInQaKC27qPMVfCHWEalhWGIs2u0b/yKvzT4RmjgtNkYIBD+xqxGxuL
YD5jb2sPHAw0mTvLwhwvmNzNZ0oD3lHSjGs/YrFVnpkwTqh2N2UlkGUQmY5bO3qI/W+cGswt38g/
FxxeKyNmUx9ROcBiWv4BA2P4xGyOhJapcCIprVVMOgkg/tzhCFsGmaM4uvQAJCdyjk0uM+5JXqV4
62sHZSss7563SbdEVtByHfTHVdHTYASeLXG7qm1BAGZ2cOY6d036TyUyix82cze+im0ZAOXO7DN6
2hvqz7S5FTGbcDleFFlVKZeeG7qVgkF6viUqiwuNWcVdpiJB6oNdyPVfVdelbUgIQlBhS1gY1MJl
8p6TRLBFysnB7E6yFpNe+gt5cAcY2r7ZrJomQWpZbEi0tGeI/t9tbWlHSM+mloZUZ85ar7wDYq4A
f48OYYvTtCHKIQDhkUB3GFqjWyyKocV8nyfb+fEh8hzrkYd9U/CrZ7JH4fAIPVpnN07hZdmO/s9G
uUyoBXgxXAkanPDmOjoPyP1XHfUGHA8NurDq/ur7nALOiGFmIIBPuobZEMQLJo5Szy/BblNKhWKt
Yu8h+rUJwob3ox86htnzP4ODxpdFQrASnil6TcsOF93DRi3915EA1K3lyXXzVVmVPD3TwBuzssyG
oj3qdy/sojNxWsnbsQMUio7owGQn/biAe44JHE/UexcKN5/wrskaGQsLKIuZAlTyWtF3tziCSLq2
PHknP4VyE4thYfGCkaafsXuV01+O7NAe1oAQuUYXVDFqQoaj1f+l1aJ/YjBfTOQgG8wtalzIO3/R
yVXThBOWlDqYJBBoI459QLqhvLPcP69ATfxKrcq5lBcrVh0E1KbrZJ3tSuFREnrMLm9zdyMW4Wuy
6sNoT+0P/JCzqFzUB9LD5WaD+lPSPShkuRyolIGpmaRW/ef+rc/jFrbQ2a4U/XYzwEXzS3BYvKwR
4PFWjhlcSCP35XyEO6/t771qvk4hNssMvI6Ed2sCuqMEoG/Df5HHGXLs/S6GbI8Q3gt03RIucWR+
K4mvuto1eQHdLZ4nxCadHDLioRmQDhGKq1WHzH03xxamiaDLg0Ky27pIcsc8rlxpxv29q2/4Va5o
RbNDFsP1XQooylpkMKbZ40QMdNPsEVFuR2E6p9Uml4IQ0u5fqYoCzC3fVRHcwdO1YRNNmAgUjT3s
Yo9jXm5ZTEkL8aigMNyyuBsqFTVuFNmUuG0H37h4mAGDk4+VN9PU60RvR8mhoYBbPzAjLSyL1CnV
8iquAwtU3j0qaqqgpnwz/EX3Facyd+wGkbrIwlODpy6Li662+NcfvhnEknCzS8x0uPOCmtba0FwL
5e9pxjTq5W7vmJbCXOY8bIpcS9XaIKfmnv6gLshhDfW46aZ9lQpqNUWSwvN4bY8tLLij5XO8Tb0h
+gGrenhhlmtmjqzKiBmnFymTSziiHdRu0eLCsXOyYkh5RFEQP5jSqDCfegv0BSUygUQxIh7UGJYL
FcqGGreBot4Q/hHcAGFnmi406FjxjjJbSigNwJUyx+5fu/M6jXy4Epm6UD3ltjeWcVmbXwG5s+dQ
9eJVS4wowboHuLPajTmAqh31DZX8Y/sAKg3/xGxOOtTFhYkqaVRKEGOgmpAxWsof90hq8/u+Bzx+
wF5/bHEL2rl4cCepvJsR57EM1xwum/SzxqZO0Iq/63lxJRuINfopfUgdthrkdyqFFO2SNsZI/zH/
Of4V88T4RF2ERDAj+9avcGlR/KjcX9cEumYCwo+j68DI75GtqAwLlEXaFo8Cc3JcYrknNbmd3eLt
fHuOUZ+4Lb/c1aWl3/Du9fhRsfsyjYeSR56Kdbv3s0JKVQzxo0Y0FuE5HVBbxq6yKAQvE1VY5eSE
KezcehgsxQTEl60eX8uCqdo4FH8Gk8KYySDCQ5trKnzMGFmTNtFy3Dfckr3mDmqVSts2eX35rjIb
bQ5/xQMBG4XGerurJU9gmRFDWVMlfmi1DRJGynRIwZxquYG00qGTiz2+7DDx1o2UWuZPU3U4CeIs
z6MHjL219NtgjTPJ2SGadrmR3krMx09p+YfwV/jCbvjdzsW3NmAjJSm6xwB2Jit3JCfSSEhGWaqX
xxYCVM8RPb3VX8mmKqRsXLiPQfI47eRkAn7lTDbJ47Voj1t9xw578EJJs214x20ctFsWimnJHvpO
UHOHdSTvQNocPkFL0ty/FO/LtVaUGVJXrwSw1LREMjwtxc2fRW08wmzM2IapQxUm+0uUDPz1UHvL
tjCm8BAJZF+NahR9kBvn/twhmvCLWEmjU47sPD+HfQRD/Z+z0JJ/xfWgP0d8/A6TxuGKnv1c4jFc
PDv+U7TJ3HGAfC6ZV9HznnOQRRjDuzgeOVUqhUr1Ih3r4i0eYJwf5xlLqEtKLiAXHBinIcPVeLqe
yNfirB47a7cs8cPnJZlF80Bg6uqxkF+Yct7wz++2wsOx7Z0R9R3GRJuFvXcTBI/9YncJXIskDSNs
JtgfUkzgvZygnwyTmx/72sMEct01DDc/cZQuckNjDcYMSXBuk/2jsOTA1fjKQE4W61aBJJqILHda
IfdQ0u6rpvCKC9F5AOB+88m35QO1ylQ7e3u6/1nMGbBZvxzVveXF4eV6Z5l2Z3S7Cmm1IK10TjMp
VPU3O/k2Fff1+9fQ4t6Om862veBSOwPaIOrgGgToqPg63+nKpv/j7IQnwiefyIAUlUCBOl3wwwsR
N6Woet3mRYIRnFGfkKai08KwPcSrYJpXwh2+g45UZ95XkxmaKlJB/k+8HBnFJwjQcV1C0LlR2Otd
Ii8EEx0YM0HgkSxaprZL5/6Zug+iIaqC5PODbD6zcplfu8TBJGm+boEVF8YmuLxsImGFzKWzaxNI
tg045HwNfHXZR/JKcpDZdP7PtqhugUkORXCMsfbW2Rbja81uogvxKYTYwofZg6IH8bhSfNVXTxtz
G/75VGqbM4Zz9dFfvErDdjiYYwlpdl6x6zchGcV6x78yYl/yADCe+6Mxmpxyf+IAB5DyawKkMcxx
iqtQOvPtDez349WbGroFfO4vpf2yrG3i+5kniNDwF6IOXo7z28TEwM763ICYt20gkLOQU31pgmO9
f2Oyo5w67YzM9NchOUxSkDAHNRxuVwEjo9r7AB+r+1AllsGWx2WQ40T2UhEWviCURav5c4qN1bNl
ywGafAtoKw72w8d2ujekcnyu2Dmo9uZfADMaTnaGrOxKv5YGDAgIbgc1DgVH6umjxCjaSXKUXi1i
j3i1rvfcxq0DU9qAraoX4A4SuBfxUy/hd1Fh66sr+T8VzkZFflsBm4qfId64bgaoIbYbtu1GkFNi
2Pa9K3HmW8uPKOBU9iVZtqNO5jVuRrNMyMvVbKzPtDSx1ETApGrSEykHIyDPgKVEn1c/zxOMyIZb
CMq+1hBZr3FqAdiBmOVQ10wqGNxey82oKDyPiOdteF+IWXHSjI8JvKVpmqav+PdKZN2mEQfkt6td
dnVR34BVYp3LeimILypo/ZQZEJYb248fMmwCQZ0sM2apEliSspRS41kLYHXMI8cFKbCnWVudJfbV
Ee7RxmERm9qhT5vhfklO2FAudt1a0hKzWKK4b8pXUHdIjyq6r2jQ+wsk3IFYtMzBQmHsuncGsQtm
fJgsF8NJQA8s3SII3/i6h5r9fMP7WEepker/l+UZj4dcS+g4YizoQWquxqd1BxNpPLs2Ll/dLQYi
DySJMitmEnLxC8wtXjZusgB5lkLw+M4xP2dIhAckIUeGSEwMZr0I+VyEdtfR8hsYcLuQxlPZRskD
ek7a6oR7BlPfS22gAWMbWi62MS8/utMlMd2nmNR4CsktoXn7dkK74/4IaoNAbLZtXJb9pSoLSUl7
+jBJLQ4Idzc8mw4xbKzNmv+beZAPrx1m9LYohnh4wLLvPJZM69G1O9s29uMsNKoXxGaFEHOCsSu5
hsPeLCsVOeuwQ0HnJjjLobyyymjJ9TIIv8EUUvw4uEggprAGP+7erw3lzn3O6KONdqVB/qr9EVq7
m9dRimUE4jBSUApIclsguvQKAl79bPmWAz6Ywa+Xwjz3dkb8VIE1Msn0oJVU07objnzExz5cIEjB
eJy/FoMW9RKDFBN05H5Xhq7jArfMwWoSBMks6+QfNM+mhQgyR0RzBPB9RGJHz18lQOXHqXzbPF6v
eHtWkeIhKjs5YT3piIA8BAj+AxbR0BkTooD5dVOylCLcHqptJS5JoYXlb7IIirSV3Q8FpxApX58R
eqVK6bfCHhinBDn2tDi7SS9pziFgqQU5WB/CZ8LQ5DE7rZ1u59si7af0Qe/HBx+SZzxz0IVUYeiR
cx+b9AnjmJUiAoQS9v5kTQAP6E0V589bUmNKUUQ+Qbxd92LH1B+mZziLGd5fBI7YRvU8Kcb/D6pu
ZKXIoM1wo3XiaCrQGQx3nrShI5drmenOxjcP95uxqLYAs+yNaSu4/P6djrbmiX2dm5D5sH+TvMIO
6Rr6P0wDY27MBJaOx9XqRiB8pBMTg5gqx3S68cRYDEE6KAdjC/8YYf+PbyJQQuZyI1o1JCrgyY8v
TlwbG/5qK9iNAFASEULSEqK51bhXWozd/jKOvvCCURo8U56oJAlwUgn2gLM8ZRSVO4tg/x6UX1v7
pf0BYHwVyyDMpiJJh4+rPp70efR2O8zQ0H0an0OtSBOCY6gdpaJvVjRzwgVYlbKtsQe0kjg6TzQB
C/f2/+t9XyZe0G/7+eh+aw0VYZk8muOpYA8K+i2kBqqyfOdxx9+Jd6Zpx2JfHYdo6Bo+GEteF3a2
y6GDzMDjHtWByZPh96rWXxgcrqylQXqbeF1pERecq11SB35nXhwFXDzE/JROq4Hy2N9O0YtUzNgy
aywgdC4pyA4gQ/w0vqmffyBehpQFCulOzjF2hQebHf/QnRHg4siv2echl9b6XhB34XEXfdmT4aGT
yy4lR5CiVnd26QleYqm7Q2sQK7evpGVva9khELrOsI/ihoVRSwSZ4iVg8njf7Px8vCd1t9hV3ykE
l0PRDNdjNEq+qMsMqv7yevIQE3puhrMeNRNZZuS5mkxI5Fmo+6OrPCWCgNzao3BkdfmzsewWaKyB
+NilvDFVyabvILh+I/4pV40uTEM0KhkGBQaglrg3rZsRY9E4nt7vwFPJ62iPC5kZQeDevHWQ33Ow
C07mllbJ80AA0632Bky5WONvu81gAd8RVrUQfuwBDU6TDa4BiDLlocNZI5r7rJQdsXevNuY6y9he
W36SFAEEF0IxZShwIr9V/G8EIZplK3H5AOXJGw75gWKqJy7nNN5VtRw3qH8E/Sh+r+LmqfwQOxFW
/7JyvqqW2mDsy3m9hoMeMwyg0CE8oW6rwdAzzwldMS4CELCU/M2HUa+cEweU+SfnPhrbRdi4kBWH
sivX58e5ll/68YlVem1WBmhu8FxNm3a3MgKD4bV8X+SbS8yl/ugfw9wxwbe9MtURZ/dSzdlUMeBv
fK1FkVWHfupIE+HvH07LbDkMn0gxswJQ3KOkWrCrjqtA64rFytPe6I80mJ+DKmYJaAHW+490ZORd
iVfG2uYDbFrg/Xii/B8ZrQk3OFPnl+plyEqjO4zOd6g9GUlfXxUoqkCoz0gE3LNUV3KWJKtYt5Zr
faEdj1eRthm7gEBIoSvLkOFsK4lCipfz5FHFaRwbVQeyaRX+AHIZIxXrsYSUpn7CPwBH8qoelsK0
80ZOEQVKlATAuSyksqgjFpyGzZOc51gs0ZuHWGs5DUhhx48nSoiRNRshMovJdkFKgFzPCLDM8eHW
NRraGqsH7jvuseHRkHHh1U07jUmTA396yAJebiORMGkqhGYIMSEgqB4AXxVCvtKZ5tspK9fWOFZ5
yW/UseWNd9745PKY1txWkY8PIj10VHs/XhEgeNY46z2ufHOHXfBEpFIHK4KyyIugidjB261Z/PY6
L9XYSxWfC2XC1WCVUcRDKvW5sgF8oksY91dnASxf0oKYsAOPb68FVtCmkQ3YNC73c1/A2aRXumQm
CYYCCvkOG5BMEHjU1tEv+8V6uRm0uKWrV0QB+YU4za6YRHK/LYfgNkh2IbhL2BJTdlxs2PJzXWC/
Kz6samUv5g3bObv2ATKlhCIDZcskX/iqe6kzdQL5B8Aws/TrBpSuw1OHn4gUqKiRLbYdFrhNECcY
U8p5SNQfkEJTgh493/l+HO9ydfI2FRGiH/XcsKWyj9/4ZTLmcyAOr8hG7GRywaKV4SI17Hwteeyw
LGI62qkxez+8w7uPQ9dm65KAFoWF54GTB7fewKVVjn7EB+HKtyE14pN345E1yk7aTlSwsCtVqGZ5
5kmvkCJaw/iFC3e08g3c7oBl/G6H44SBveAuzkvII8gKO1kHty2de/AoFvPmrfL3u0yMT28CdZxl
W9RuTDX2ZWiwXHSrYDkhWWHzlnv+EEdK/7tbB2whjUeRcXuew9iRU2ygTmo/wJBnuWDMIxcm1Y0Z
8YLQrT3qneTvgbRjWu0YaSLla/LOhQdiF924fwkb7lWAsgWo4m54vAiYJzkmvnxwpt/M0bIVjBR8
9ja9XHq+iEvBBmjbgvZVygq1s3P3HkP00MB5uRYkt3pdPGVAVLPI0fzf1Blaj7GokhSHv7iH9hk/
CmMhwBAETE5fT1FNxAp+YCXTyzxG6HZNOXEm+AHtXfAxUUHvDpMWqD1GwGcW4FgNfM88dsnVEH8r
CcwBcqhC6TqFFpJTybmA4RBCpllxgW88ymIExHmPfSUv/f5JvCA848hvJBDtaGfoWRVec4CDd5Ry
y+7G6n5MkP8GtjXaKqUmH6cRMjILvb+4yBriyKb74A7VsBr/J+O8zu1cf5ful9wT5kdaJGdlGpcZ
lFDYvDN9A+N1FTr8xQKFUbTxGoOqS5tCDm2u2YYKGOnQueffVHmV91yWtNO59W9SqJuGDvJ/3QeQ
taGg9SRyKjvjGGyN4zKSdykAY7K1dVWNcClrpOYKbkiMQ6ONDEaXgRJTQT7z7AJ9oSes5L5l4XrV
2ee8yI2Lkdf+64n2LBOgWmkj0M91LcGSN23DzxdSm3zEW+OOeW6NlOrjZQsrLeR6amQIomXsf7sX
aFXasP+UGvIdgAPuL8N9d6rzb1pWVFW/0MYpzC706MKxxYLKpiY7Vh7PaJdcac3ddD0+IgQztJVj
E2NSv9U/TKuHuhsR+6fi5a6pdzKn+20Bib3My87bkjztfxBcZqQHtVDodBaK+W2o/w6sBo053s2E
cF/axQVXsWjpjma24A21Q4kAV8ktPTZgT6iFED0sCD536l2HaPs3dhwqllr9a1HnYG6eN0en423h
r6Eg+0U3DbC3ZX4RNwxKeI6wviZOVzFT1Rqe1jmzOtO8nkbB+kxeEw9p0VoZpv4dxpgXllTEfIQF
99NyZmdPyT26j4eK6Reuu8DCvd2tiK7nN4l7Vtfnz/o7x3nhUW2PMMV8BKjBLGigVa0it93yXWaq
U7eXlMPdNKKTobBC0zgOR085xvXxwY7qsLEatHBzYtQeDsGUP+SE4SOmSY43epnaHGIar3Yi0w41
K5n/GADv4EgJnlvO9vwwfjDOEX20CyuO8lO+uA1ggWX87o/QL739lxxtmnjku/R9L3UWVAQwl3TC
3B49NtvNcTJqG1L/aBeuXLa8DI+UlfLfCr1ezISCkiF6QoKIoG+oPAuxD3h9asjHd3nmBzq3ySQt
bZNBma+l3QtIz3NgunvFyvrHJMisKpH0xP24CK1/HU8ZDNPmkdLEDrpZSK7+UuVbFaC0UGwtr8EN
Q88MZdpLvKSwWQyBRmLX33vRFM7CnNuZcejbw2Y3IZvtS+ZRlwMh4eQ+dmaQ0yovS2GPQxn32R4D
sNZZ4tIYowRLk3Qoc6FijVNPSdX1A6icsmWalkAxUU2XjXq6IEE6E7vBz9wKflQMj6tMiFtd7Py+
2EnHmvsCHEgE5sDlcN1BC1WW3kX3yiL04I+rnvcEtxquILYsZQcfU6M0Jy1FIQHkq3rPkhCA6V6J
fD2MHZm6T2vSzvkUGVTIMjLWZLQ/ew68QwJLglE5rRnI91eocEJkYmzt17YIpQQu0f51lh49FwmT
Aev8ZQeOMWvB8rIgf/WDB5ytpY6/UX2TuNj4ozNIfBmI+xsiInd4iWA5sC3OvQoq8ABvBEUC4aYJ
SYqpu1BezjeznAf/X4Q69hsOfP8fy+3jiAjtsSz/QCr8xWUcwpMGSSo+QXHN8WeiBGJBZZ3vJCFY
8XGKBdmqNdnEriFGAx4uSEKtRuxVWuJG/1Q1GmlE0Yfge3SswiXo9Jf08UMXheU+4/Ulkio9UrSP
oqp23rejllJfXZ4AZjFaqIvQz6TUR8yjR4TOgNUXH7DzjHepJ+cSKjO9lHViQH+rHq/Ck6WuGcJw
1GnO3wBtTg+QheHjLECUzJGq1P09DYsSooryg4Q/GTWT+cCRNIr1gTB6G3bc8kX37G12jJAo2gb0
4FLVTGuQGuj/7nluP5fc8L+Z3fIqNdkzo0r0XPn7yvDRufacZ6HvspxG/Rt+hr47hpK0Es8Vj2RM
0B6rAmdNsCVYk8QdlSLvxlU1EFRT1h80+64qeJDlKfpHk+3H3V7d70fEc09QdEGJf3gXSTkOMGXP
Ox7KO5RWmlLVEihaDa4YePVevLBCVkWvZiEdpj/OrZjjaQE3ybMJ2FPUG/MI0X1owtpkyqB+SCJg
wh+IWsTJ91NUtWMG50jTZoPN1k/w0GA+9bjBkE62L5tzTcHyhCClKLiXry1BpEOUhe7FuSkMgVmC
4g6ilF/71rFV4hPE4YXHYBxmlMiyFuGm3sdZEMZZ+GW5bsJVf96XY5vbAQ8YLCDgWML0km3YHKCE
A4OlBKP1NZDqQ7hFNUKcBWfmmAF7Pm1BG1COwDpMgQeTePXVBX0YLKpoQPfw+eHwPsj2e3giVqKm
Ahsd9z6K6/aSj5kiBQyUUa9nGnnRNOtFf8LEsAulhi1y3rNExIwyMkTBepLLKGSmLoXlLWzsTFIl
4QCmuHYf9NluVeSz5+KZzLuivUP3/h27WnjBH5Q4te4E88f+9mNKTPxtGuOR5CgwXi2Rb6IpIJ0j
Sq5BYOMlGqFOs7sKVjYgG7t8qmeu4NYfMOT3G/bJOHMEeHCLI9t35OM1b9vHDt5zRATD1oNGXUpm
4bVpb05GFRtm9VpB0TD/u5GaUrK58N000b9Fc+IFYqz/JXAF4JxI1AgnQHahyCvnr7eV923BtsCt
XIB6XWMTUrmyPF45gzzDUvO0Q5tDJAh/IodvJ+y+uSv/iaNMhQX4fVDEsBztOOyc6FDOdtFYkc78
WI12gyflXEO52pLk3ixguLRP7cyOV0kflq+uv712inbdlBh88h86pgwTEQZBxhZqV0uNXYascYh3
ppXnmCPDU10uiQk3U2Ey6CpICmLy0y/ca7+T2QDMUyXFX9N6n7IFB2oconqkeitl/bFQ+I3Fa5wo
SnEClE/7cWGXkW6W6Wj95P70RKuhX24e6asnVPdNAWW3x+PQwPuQZzMNBHbzhVUzql6zEjn3HyHj
v2V5nRlPBKVKs9uDO2LXN1Bx2xjWePk8FNr4DM32E4EC+FjFTazq7HuT34JX/s+z2f++oWxqDZ4U
1uD5OYOk2ROjvexCjtGNU3Q0WoSypC7dasSAv2Am52NYf3QoYlz8682ZzW38K29hT9MKnsITPgMT
d9SM1Cj/L4I5wo42JbLglgxHKy9ps4VDlfHC+JoKcQXphqLK2LJUmiW8xGod/fBrAMQHX6sWA0HT
/V8FSulYPsR2PgA9CWAQYscDey76V9VCDlLz/Nz4SElHUoaQmF1/1ZYOSmhYsdhpvFtdHeSX1QiF
j+J6g8QhAB71wVR81/natwwGOvmeDDgiATjhdu1sy/Sc52fD2iPDK7+3BNfxwq4itPtYJ8TdSYjn
rODkdnm5udNmWVROnZ08kQ9gZKsREbx/evVvtspdGe0WKcJWC0xesZc2R0s6V3JcAthlL2iuPWM9
LXaI5IOL3VB5FoVXxSj5nol9I+7+XNxqAC55P4IWiaBE5ZyXmVkXiNvO+uK6X+6xncsWG7Cn3N1/
abbhxg/GKa6YIQx+x1SYonL9HueSslsqucXr2iU2/JkDKmwUmzUcwooKIKGmE64p5WOOZHpAeTwB
p4eMbruvycU57Fd9nKKP7/z3DNG2w8XZlt3px+NOCEAhRH8NGcx64U+ail7WU2asyYEkJ+XAjGRQ
OskTU5QaSA+2T016pmbvZXw0l3ITBV67lP5oylydMO/9FH1p6skyuNnJjsVvt9fikypsTqPeJdS2
GPZoc9j8S1JsOtIGivokg0Z5nX/NUDJGpPG76JXx9GdyR0M9D7InbcAlnFtyiBrNv0vEN1okJVv3
h+aNurfzITSoIV0aFt740bZkN28AxqmptLdY6Sh9LPfycvW+nO7NeHGY53lvfItXmbTT9gd7efwR
/AdvG7iRqHMlVjCHCsTfzq1vXxCZ8ecAU75YRcxSUIEdUAtYGUGpBfLCUEoLCZP5qS5V7033xOHS
csTBP8r5MwI+QMOkmS0DNPrxw+DDaTJJ8BT6IvAPRC4PlcYZBLrM+hRW0spseyGqaRtr9+5FpsAZ
PBQQXnHkiHvZfW1sedy1ibiAzxy+D4qkxaw7sLzvBC30NJnmVx3LF4oyTYnh1xGnZGpbuTE+vCoM
8zP2o/NKya2K12/rlSmbiGvwjugOJHwrWHzIeojryjMkAGyUChA7xBFImgfbXcpExeALeZlZFz8W
L3yKvW4uKqIMQ5wFrM93gXIjSRtFIPRDrJJ8HjdfJROSqzebiSxkmzzkc/1MTzd06v84nz+1Y+2j
PPdmCnS7rL1uHnTCk/vkp6jKIHXuS9whzn8qENoZeViLi8FmYqLMVbbB+J1F04A3yEP8QS5b3gtV
elNH7gxZaf93++Wq+A8VBxUR94ZmxujKiLBhc5ShAOpgTDkXIXlv2bTmKX9WmItr2S8Aody2NKuj
ALjtxUa7/rMaNwmTG060Ah+9MZjFjz5exZCAFzZMD3YSEGGQPcSoWC0TDUf28KHiMphCcK4krLhy
le4K5LCaTUhsUvaJCzmrOhbyU+EK56ebNXBufdeDQ8BE+xFr3XROlKB7aQVUKfoDBppPpFADWSBh
DvVMfzOeVk3qfGopPa7CKl4rieWfW/QiFcw2v0H915d9xa/R8WRHEn7iKUO+E8qT97RI21BkCSLf
st3lbyJgR9fPIfU8CdtCKMxDd8fyUMxNKav1vctc3Au9fVZGQfN7uOiS3JbG37GKZ+NquXXT2uzQ
+9BogNBPNkkmp0akWsIf5ywxLb+IPE2Kk3kGIoVW4RqApyXS/Ez1KRFApQ3EKyd1sGeUknpUXwMd
aybfKOsPgPDBIpRiNyVFiNqs43soLUQw7ce5XgJelVS+RMwISqiyB33MvZbojAfJnd0tIZv95kv5
wv1gzkdEZFxXA022uSo3xy5RGOKa/poGZP8WElM4MJzR1mSbr0rdNyqyBDwmv8/tDx/t0aQc1Vzl
MoyA/vWGvZ/JKSettZBGnCjiR4j3r8LygSig38FmxL4NejJfQSwK2RzWrXxeeet/ifff6wDAwopG
9BaVXbIZqpnMJLbx6Jrf5Kc9++waEn5OVQJRkPgiQWIPjDfLzJI+/Je2tr8TaQ1F2KfVHn4q0Yii
+JeYKzGSgPQPVzcv2UeR5R50AW46JM40JOHpaVjHA2hJpDIIgLrvtEVjhe6F8UBayZHjwnJmp2TJ
OD/Cx2jzh0Mm0K2UKhgjbXCrI6B8po3pr7fPXyKzJSsRiI/ZTiD9eUW3MUHcrgV4D9cfxy0GtLDK
UYz1Jo2NrI9xrC2g/ebURLh2cqtM9AbmRr5HyT2rt1UUHAwvsuY6aBfqLluOyw+dLJD9gqsfrDZA
h97xt/ouqzD9FPBqJjOaGjZUGm54IEdG5sMkoHGaR+4T7nYROsLqNMY/Q/+tRtEdlFonc5l883LW
vA4/BfV9DlV0eiLwwFs1VdTlK2MOSYc/wqYZoV/4Y+PqB3h6xzDy9C4IXN4BF/xED4Huop4DfngO
MuuodPr/mv1kknlfHgW51VN+R3ZkTsxZmS6FIyxW2tNeMeGrN7Z22S+sdk1IKhOtNMNRWIbj2ULf
8eErAu9aVRz+9MPWFpAB+Mk5DUUSZ11y+Sl24d5e5eQ5pdEiqWiP4ZWWJ1RcuhoCGe6vUEZEuaHB
fzUQsA4Tucdglxlue0WmPu1n3BCbaGj5byqzTourdk0xXFyvg5/cUfs30xojUFSBs9tdqPPo19MI
54k6JiyU7bE9J4mVqyU7Tx2dcBc2kyRxGyvJizANqIEP37Yg/vCR6dIc1soOm1LXKTrO8twh6gmv
lid1J/Nsxe41QPmFGvj5mUZifmEqq/oi1UZ9DN2G4ptTLv5q30N3a2V/B9mLeDCMOxNRdcOfa+LG
LUrfXY8H+e2qh6Do5sodLjyyfn+tkSCgDrL/961RYXvUBQkdH2PEp2PD4KSeO9rEn6eZMqnQK+uR
lCB1jL7U4mQfETugJ4Z1Jp8bQeOh8s4JcRs+aEGMl+AIUvig0zNluZ3zKacm901+lG19wv0xThNJ
0j+NNg/MR5oUm5aeNlLwKFDBu13AzHUab1jVA8pA6Z2SlDYik8ZXAwYG6g2kdesBU2iiHKFbn0z+
3IYyzg6EXrlJjtH8VczVqYPhPqcio5mbJcDwFNSv4Id7v28GOyUZ66aS2IdCLLP0bdFMskd9Eon3
qPTA8HV3oOnKQSpbfQVSq1OShf1Ei36y/QI8C/LsNd83Qr9vwpaa60XjkVHgP6IsKxC3C/VGBGUe
1e7+6HZs0HQlTSQBZNIN/34tHf1mCwQtkmdHwvr3/m/jSYq/SndIcnSTb0fi/TOTicAeiIEs8GI2
kc82cV2DYNELH09BpAmJRxBHGumE6YTSk74yP7DalfL0VKxU4HRgbQnOA9Dixf934n0OHKRcKAbH
rlFDll2kSqsLz50HC1Iunlkbt/kDkfR0nvM59RbhHTrLYLLJfu1bOjHo2L/53fSDKIqgl54fyxoh
Qcen013rk22S1yYNEF2IJAi59UK6H26iCAkTtAZIsqfBvAPBqcqorcQSvlpuqGR7v4ElSQDyqugM
JyZfaamLnr91LrAQFfpM7LUioL1lRdNH8g3o7jSpQsUlLhNm/q64GaPbxozK/ky5PmmqhfZzryc5
10Qsy8D4/FzbR0bC+6IZWpc+svvxg4S+9JFLLV1lpgzhVIm1IdbF+6rXf1+x++RuKUiHHuOk8png
H+ogEgmlg8kZfrZyNNG9mDRnqigRrI5bnDQ331hjY04xnLpcsc1ad2g8PjxbMKEsghvp8OwYOBIY
lhNXZDt09tSPL/N66TeFHFUo2rFevxPH5SvLfG4L5YAAI3RR5RoTWSJkzzqCdNLO+dw0KRMCoiNa
KwvHYOqMUwuAxgN20E0QmZV5dYSJZTiQ1pRryw+JVPRWukHe4WeLxecCo7Qyou+LZtoGzOY4yqhe
LhlRSG6LOE93DwYg122KPggQLX95izmLaIdqGMmkVoxuiG72k43PYQADDJ9+3C+rwfG4q2qwQEXq
vyhSdF8RWZzUwaBAzNEHt9TWJzUbSOmTdhgxAcvaE/CghejXJ2jcmDDuJMqt6yZ5GBf8dnqAeoVJ
WBLr2jnT3uyZx00El+eNEEw6vQFxsbH/NXEOJHwuWV0SVBD09ul7z9oPfT0R9ph6zVWpkBlwcu/F
BUpbMI72daXMKZ4jsG5LjSDNtt0fHV4TOqPqObxVtAZ34ibHqChudsGymJ7RQ/seMeiT74RDMaCR
ynDGoqnlT8zIvk/Bgs9CnqkRCrfW4HFfNqlOxZKPGu/x1EhudhZFs5XL1lKqvs8Xm04YJv8vQLZt
GOp5LAcOdD/u2G2Vx2rr/qML2lGQzEYmJFZOx0t0ap+DwiVBtICqNgdUpCrB+rmHAIwWRMyXB0CR
wl0DOF0IlOZ/nBjSqD5dCFVquZeenoeSJN2JRRU/Tu5p7ZOvRHtxRrLQx1D/2WkaHASF5R66KrsA
B26p4PRwrRXQyMUaeohnJ7zERsAS7w2+aizkzQHfwJLvgY2TU71CJSX5rLshtlIvAohvl+VirA59
Nbgd0LQxra8qE8VXhLxkVNlh/2NNYPZDP/jMVX706YpmUP1P21POiRNfRFXRcGT8c5kWlEw4d7ui
nJRFtwXenrBV1wE/g0Kxi/spxmsk65rv8TT1tIEI8v3CNEq0gQmjtJxSPCJcu6qpqpAc4BTWS7xH
EAywmfDvSbG8HpyVwP6gVJK4NiVdJlofbMwZivIY0S99aDDFHk6f3N1Ezpf3cmdWd84uKh4PuqHI
gL/Zaj/OhVEe9I1/8m6WILl01kpDTnWyuPYSWYL1T4qIYuKo8EOwmbAYAtNRRRvn3G196iZ9BY14
zSAdUi/1x3vR3wwb1J8UMdI0DvnWAa8KLYMO2JpBAh6UtkxCFAoeBkgVdawGE28njKJKA5IbkzeE
vMdvyt47Gz8RyajpkdV584YzZ33mGUByCFjoDzhPi0RPAat5YZKmEBG4ClY1q123OfbVTsKhWVf3
+Bu6m2HSEJr978uDfeXUgIRoEbJu5lLF40mbIuwFWZN0EpiXyuuCWwUsGpZgBcX6h0Q5MrJsqkcp
etFjSj/mzH7YdoL0nXKLbpCd1bIdOvTRMtAZaxRpD67TKJ5JKGTayAK4alZeI5qkt7Q/e+W2FMMk
YyMVOpW9hhjECiNOI/J8zIa9SZxoLo6NQGLXNRdpBnsyeuItxWWMAXtJ2OJfK2IWIzz2XW5NPF7z
DGaGpg+bBhVG4HawdQiib8VhLMhOVQ/MiGaOtekcjzFgr6ca31yxSl3HOeSth8RIOdYUT78106kr
i+gqhSrnXpqP3KT4Re5ZCPDSSo9LZbRFEdojGfMxHdtaeFEHcY3Ww8moST5IyaBkgqGOMOQIHUmR
Ymt5U4KxhoDPSkKfYrLZV3BimXVvNHevCKirxFzQGuNNXkXEEf+TBQkTYBMtsiIS+tR3K5uMqqVB
aNETASaAAwaRw3//NqYWwwyBX9vRnR7dRHi0NCTivTZtIPQ0v/dl/FF1/jGVq+tlWMRn5BKMWi27
1FBeH0DGm94QaRTxuJ62xr2ApVygP/+B2HUvCCwISAkz9A5LVd8nAlr4dqPrXYTJB2xTdYbxHXTi
ntRcimLhP7pR66wemFnVCxnPFuJWtgkfThOr4+JXQ7QYsILqEfqMhg6db3pXmLt1zT0J2LUAJPYw
pzN5/4Z9T/brDFh50DMNYvovdAKaV5UgxPQTEghkL6InY7ysAglQyvps2gPMrTneHYbG/fL0J+b0
47d8gh/8TVJkL/+opqebfQkc8oUkfUEP/sJxp2vycGSJwSK4VoUQgVKeZL4WeChyr9d85hbmL0d7
dRCtvOSEE0SBFuT9DoM8G/rnD2t5yXFaLEIDFSYfP3JuUuktWezfLBPWVkx6yY88PVNPW66qYEsu
obbCXWxxoPSP3z+UyCzKaRfvQbOx/Pi0GlyF3XbBzp5vvQmW3m3A5g+Hm1P/7gw4sfpZa6HCgPbl
Ox9tfUgb1pl4V4idBOby5zs7OMIVmG3GNASZXeXZfl/abvt5gacO6U549AEKEZR/yDTDT3ZhW8Qg
qTozuUwfdvD29g1ePkLOgtQyHvocY/EMCAUfMfGGLURu58AWrtmLkbbX83Z03EMJAzqSeBdUGa24
QB0UgY7NmYi0QD+k0wNSLxWyaGTmAHXL1r7X8sH3WbTCWRnYG51O6mDCJhtR+JhQTO1xLFLaIF2D
vEiGx5JTjcqL+91eqCJvPnmLQjw1i8ai00MbCqlEXS13uqp7y5PriX6kmekV1ns308VUviTiS0c4
OUOIxKIlkJP4KQ4LmwMuEKw35cvHtlDmUzk3KzHAIBtFEinCME2G2YygEmC+H/yev/gnOBUk2sJD
+i0jpSktUs5iCpzmJLXn3V2NB7Jri3INubUuyTOVqEufAHtK/479nYl1tbeI/JzV3RJJHX3HJSpp
Z96EcthhwItXuSajCaqZF+l0gwqFBLy0lBJlj1kCw3BTlgMECblaMrw8g2stJG0hXz0mCkTMnM3L
1ngnkgmsQgcnNANKAe3F/qAgL728ZUsaenpQeTgzAC6QYPpY806LOYpvf3hL+i7ze90jW6kwN2rj
PlJmGpD+4u5cG389J6a0h68g+w1a8RTxFn0T4/SdZvw7CjCAbPJAapm6x81/zgeVW3ylLyyxVb+p
CEVGeYcRLwJPPnWda9owHyu6WeiAePbv/b5yoP6G8JSSVBfVrW7Ct90BX5MtNPuFSj2uC7HcZlE6
5KS91Q43tjbn4ke1jM/Aj9oYM6fvdg35+6NUx42nDfxW33jd2MI5d2vqPUTv8O9GBEjrhx9gKjmh
giZYNqA4CCpevTmDIx6+eZrEuiwpUN7chW4x7vC2ssZcJ8BFr+TUPH1iaGsNSYcPFoBfKZf/beMr
KYMZ66IAVXHBHlED+wIMwm6w5Rjv2BUImS3bp9E37Xmu7Cn5M0istTNePaUOA/n0k6eHdLGZZnGN
cFmFbqNNRtGMYpeBUBWvPj/ndymQVqP4YqGgNv6NI2C0Gq06qk9YUXCMJeXXEKKAFq1YhqKzA4JE
P6Z8KIQHQtamqFvAqurAmug84ReXrO7gilKEzEBs1pD0Ta2K8p1nhiF84Eh0gepfXxl8yxmwXozC
dqb5vtcYHtzmEHt9fpxwS2vjwadB1lWQk/K9LbROmHzHdZmM8TOcWX9U34A4zpLaissX4rCYl/LD
wavg/p8WovEM3Wh79qgRotg2Hkou4T6niaS5ZAwFkA9WXPc24TmMvrDZ+x2uPfikh8Hs8W64KtaX
Sf/RrLRQ1ZnXC9374Ssv2el7vMYoPRAxQ9Bpf0Jr2ZOuNeMx8Vwpvd9crT2qHHmBrE1NE1PwzK0D
NOB7i45UVOPEmIUn4NcBE4mvZVybKKEyGQnkBVR0q0npmknrURJyXdlIiELbP4h3kb6FgWkUjLuv
dCM4Ohz0a5x7wePrAuDAh8dlZ2/6tIZembpeVIBdbjloE3dUXFS6lPzHJ1xHsmJ7OAPtCpsxUJq3
wdTWxOljmzbGLoMUg2/E7kcNX8eT0eWBCeNqdg+PkQssCy6BQpswK7hyFKznZw5YCiRXVpNH3MLX
wJmI/FzEZ4qt/EtcLSHrYt6DUKDP9GwH863IqbIqjKCbzk1GtkmvSqleGcCtva7Amf41WavgPr73
+GeRvzhvofR8srx4qNm/I2UFqhGhVuLnYdVoz8ct9Zo+1xNWNGr5JjWNHYdhR0eekcyp66gZHAB+
mFd7CQz6MLsbKHwmueqwubxMy7EY1/acCsx4OYSIp4Ru6aZq+OxyeKRUXliRIlRATUDbU3vKb+x0
EWGAKki81jetTA6u8CF+DUrgY7NRh6XLqh+DKRXWVKtbX9PD1DekPgOQEVevZo6KE3XSxuQpR1E6
BJQqip2odW4dp9woiOb1IPN4AQUQGFpASOgw0c+uOh7RyKrsXiTwjvRD89ES9OQm8OHjwqzuX++W
dOY/aLYhN/w9+iw4DfpZbEBsRyrz+hwYqoYQqxxLYn79+TpdzMlSyRFMlVgy3m+gqVD071O4kr4J
fcs+Bdy7kPbdAO1CjRvzs2UUL3US7uoUdpuxnw1DgqhbXVDvgBWa4nSPtbqPR+5pdB0K9sjKWtGY
1jIv5Rn0aTvcE3SM0De3+Se3dLRrXzZak/APbTYshDi5/PEvkDgUKxtSZmld6ONTJ47eNwtKt5r6
IG2WkGUrXfsquW/UAl9gWT7rDNw3O3/OW+ULunQDPIF0NQLXlertkMtbYZ6djxj0p+mZ3SwddvT0
NWqVwpdiUH8iaSoUuMAfYWNgYydbR8N12K1SXhk4ynzxBINDg6vTCilqkENskg0vPS/Y3egSg89s
mTIZqQAAlO2sm017UIgH1Z+Uv6i6pqpHxxr9UG80q0lF3cNA8R8bCl0icZvsVO/DKKsOjJ5N7iTk
B/1oiggw5eHUXSgwD7GfrsJ1eIM9tmIE7uMrrhARNl1ArSyb1BlxgkcjjlW0vkMBemzClNExhcwD
SCT3YuqOryRWi+/8lcCMi9kZZg5jmezw2TABW3E5gMOjQzgYSi+ZryeAx4BF1JOQaz01woPjls57
BqZj1teatCs0OIso2h5/MN2GMNW3prUtSftTKcmOQ75/mJW/XI9eQZa0nrgTZ92xEFD7hy/TVdbq
M73BWlvoHquS5AMirSaYmShT68Cz/89MIaIaEqTQ8v+nZTTdJLD0u5biaNs3bsM9jeX6PhZ+LEFM
Ry+2OkJy+G2z21081GNViGu7uW4yg/93AAkLR4m1gK+BjeVyDjkwWIMSzvm3UVNh5x9CpFfvsgVZ
pzfHu9StymecQq71BhULlmjBJ8gjzRZ0uOfNTB2BfPofT2F4/a5HmbWxzWsHMjkaIp4lQvC0JVhV
CUB+syX7ZWytbgFlYY1I56ztZ0OU0878K1kARZz4OCeaIGwbilW1kQ3+yhs3VJwJqnFCWvRpPDud
Gm7SOjgbXt2uh6DFXX6NSQBZtEim8z9yKNXZ706AHG2J0hIEZ/DhtSm/Urvz00Px8vNfaVfneiN5
5/bjk7Q8y+GBUP1Y39kTsacEWpv4RD430kyfLSuRnJ1dXAzVm55Dz7B79iwE49Xi2XzrLZCCiFBr
a095Z8WzPphaQ/lR4CjWd8vfxQATBvlmXBcZq6xaW4wF2UgACOHLUDyWDmP8eWAIumD3fWDiawav
uVz78Dtvk540j7C9qth/w4FC9MIZLGVQiSvlKK6Zv8d1sVnW7lMeXTF5IyaWa431P/wXMj8Pk1tC
2thGEKNb0nON2gUi/Qq8o0s63K7eTf4holdAFUN2e1SfjZKP9HU+Dnj0+zSa9bR/Qs7s+Q5Qzs30
plbq4c+WY1nwjd/a+4c9WPGFWNOzf4LBGQyrSE6exN0h5GmahtW5vn0r8mf45bkH5RKXIolPuDhh
+Q7k+waNjgAac7Zp5Izl8Kv5pj3VV21WEebzFpzsUIys95xSChDrmXn3pzL7sf0DfFR4xQxMeK9T
owt4kSMMERkjnhcZOO9shyEenys9v07EsnG0AlDN+MSFvcYr0eWX20C3Fbe4C7PpgWDQu2xJBBAi
AP7hg+b4N7cFKrWchBnUDmuz8Rzu4XHcn1QnKvpw7hEN0PgDYPzWy+rqgxgmaQJbkkFwOYxbFBGR
tp3LTvcZRaOgL0uglRe1BqeWH0wumWWkRvosYyvAztSoLoiGF9gyw/eLsi6lzR1wb7mIPGDiyCl/
H2tCxjoJ9oi78hhKeqU859Sf68QjioHiYw9oowfJ05SyKR3rv6oGV2GrmR0vEdyrSuXuCyLZCBdt
wY710RAlyzpGJpvQQF5nCQ9Jrks4FcuvRyw1PbNPQCWKTWaVPkNYFwbg06f5J9toeNMpMv07U7X0
T9anrJwL4ZfhM7ERsp9wQMJ0iRUZ/DJTl2vFDvICjmmom4MaRCw0ZJujkIHfAKu/GnQGtacArVvk
e/1abHSiq7UcraeeuYuO55+3EfSrUHTZFLfB5JNXVL6sjcXhrF8IK1oHxheAvWh8757YLcoixsGt
fkFtxTMwNnumkWeEBUXKs7pK1NkQuNbNhSziAou+9ElP9Eisf+wAotWDcIE4dSbGkDeNrXXu0Pp9
ZwBPCa/gwJxMlyJGBk1yolpP/eS5Dd6F/SJ3NGo4l/Yd646w1mlZoPiO8ziM7y9pcTQIL/sWPGIQ
ZXjA7SKECB+sVrwDrpPFqe0G+Y2V0SjRIXaF/Xhqoa93huUbQIubohdOKw38b238YEiXG9ySq0/F
x3DPVWVcDu5vilFNhJoe5EJmSFxDahkF0yo18Qmb55RNdH7yiU32UYRqRS+y+wtjUAy+eZW/TH+Q
b9gY2/x84nB9t2fjWTX2NoUOZK066fHlKlVcJsIfHy9JP8RzNYxjeg7Gxetq+Z2/Y8w8Cq5j/hRE
dgCtj6tPgEG5nsPwLVWsugvtdGdyI/xNdg7pxfxZT1+AqHTbeQrNirOYFXrZllFPy4EaIreU8rtu
sJVGSsoCS7l7/8t/tEGJSU20eR8RrZ89pGoIgcXOIQIR69c1ZpGTvr/Me82lQ2gYY94jDjtFOboh
+ceYudHRLBfUcH71WbRIq3WoNtmTr0xA4uUK4eFoBh8NUnxyy8V6yUMqjB1jEFuhJb7Zxw/ZWjwm
aTV6Rgjm6ll0+X7lFNdWScWemUEqPoKSdoj38ZsL4eQgUIlM0ubzwCCJf6Dcr7Nm11rsdpiFPnA1
t3A+QMoqgFDFsTin7nfA5w/8PUUK2uI18XUhZJvndU7CWDuNGFG8SdVT7Rnvve/4sXBH4IIL0IE7
px/JQn7KJxsGxHL5wHkmd8TIQagX+I5C0UB4x3Z+61tEhYvClDX7o3nnu+L9WWK0MpZIiHbbDE6D
j2hC2LvS361vDrD7hEtgtI5MJDa4GmyJFGRyNpTm956J8o4o6+Dx/Yy+6Xub+NPp5svN+7J0Hy4/
fixMMihDl1Ax7WOJ/+DU/+zYNWk+Rj44/rOzGYUf9oDu7I10kuBxuygzIJAwLpU5FM7ZdehrT19y
wjk19f/DpCFyOAmdCCSxIFbsZIW9KiCjiSR31jKWkaCHSDm+VGa0T8VgwWvNvBE0TnH2F4GN/NSR
Crvuw8Rk9BATO9kCaHkScnTIQipamEYLCcrXtBebDKfkg5z3mzyhOugRgHtIcW5e5J/tZh7vlgVh
J0VW5zQXydrMYm/iq1/QECupS0DBQTpEKvSwvNxBhVUizCeV4DxzKj7abdVcLnqgY/YkwtseWiwW
XboAk5atUNjRISr3AyHtlGc4+PP/+mYRaxDDw+Lq+Q3tsy/uNN+Zg6hJfNmPRZYasBJ/LHYgB4uj
zOarLTULHFgR5gTx1rdmM2i+tuo7ULFEXkN2pKkUrWKTjPo8ImATmeBukVomHP7rYHT81KXxu0VV
NtVnpnv39nzm7/cqXWWSf3ChKNlgKaONc4v39QuEscKlQj7mNTfcAcSi/60iUH5ZRoBugsnvIrdv
X9jPuppSIlOoHJjTiKvM/rapTp3YYHBfJ8KAb1wJiF7jElgWGhSYn8S2Pye4IuZ+q+rpaHImp4JB
5wht8Pd9QqNPHThB5d0B0HuT9xQlwkwIXwWn8EoE1FCdlO80aVegM+sjry03RLs07K5n9NQxn06x
FKv6jmffQA1Unbzx1CLcu6aD9+sTLrr8x77rpy5Hoq2Q6UNf6SUGy3DE1PgzG/rV8KZfTKbl8/nY
CBMhhVNXhX69ClrBmCHWG2wz+RhkZiX+YCMqs5sn8eMkTyPZE0XGRcMqPWtAax4MUZXqXoAtWLpY
ca3j1MIKi9JZxqBPZyCARnFORPFBM2t6JTzofehcYDw6BaQj6ugqRlim+AdA2QwWKGrXWBmQfavj
JuEAw8G8aNc4WhzW3HkwSWHipH2BDiY9nainxY6rZTUTg0JzsbXPEBMQvXI0d+LN5Tu1Xg3x1Cul
fP6yCaWBsZzt9yLp4ZCoPVvj2tyqmt3pBZmyXYr4bRj1Jye+qhssaolbnaA1ZPH1MJJBZCxrhgU/
/OnRFh1att8jgcX4jLm6ap+5j0hX+pxiH9HT4RIazStxcKxe0kokwjQ0Gizo4UCIpD5W+c8fr0Iq
Nyy9MUnwktVUQdnzl1uiVrrWgrZ1JQUoiKcOJc+eKbDGlysEZziytHftHEtAxExNyboeb36+Y9YZ
Cvjq6NNZlXqnabYMTicj/9yt76l9beX1ZFc/gKto6nOOmO/VW2NzRo5uHFwj3fgTnnHR6F4XWttU
JEafpyGalUaQJGUnoWCBiNZkdrVZwnCPCr9hVcZ3/VmdTbEX9JsdTM3tEH3EE8w6BvsjeVQvRFjp
LwNSwfKGTXZZEZOvaagxl57a7knmir1pxEnexoN1lAnL/rWxkCjDQRnPNNXSUWJGGzVqm4V+SzNa
rvVro3FE5p8przkkJVbExuPJiWy4cIJVGKbdH0W79KYyG1WhjAFi2mxrUtSfq70nIu96cmFzF2GL
pPPVF1JmGNnfS/iKE+0XHB45g9e2Ik+8WQV7EKlSEKWyrD+eqaJGwQvQSKNKIv8YbJKfV1/gBegG
XBNJqlIc1gAmQrYzZTgF9VozkNoHPiGtjd4fsM3DiKhXxKZX3Ed+efYHP/PjQq8W5EEM2vSGrqHc
jWzovkO6AeKr5/2U2/7ne/zwtovpoKJB8a0HF4o05dlRnEwPqwUBhDC+h4K+jVBesP2akijLYDV+
eOdOKHqbfVwiIICn7kjV5+MrvA7Dn86rsgGAwsRgqM6IZg2yDOjSGrrgClo8d/Lod8zSm2exYgYu
XaSg/U3ZkWfdrKByoKutvpvEL9sm64HWJef5R8RUPYU8yllmRdKmn+om1vrihx2HxUpwJPyv6JtI
URTa0CIfsbtpGMEooMU0QkC1HInGOf5ff506HuJ15OSlNeUPflUdcgTWM6Z8poZHZ1pGMZQdfvhN
6nrrntNPwZyiTyEN5vc5wfvSFe45871aJUNhSmtx2ua0XsUPVx/oVFr5O33UJa+qbk+uMBQqOBXf
/TprTVZVEumPnah6yuLdPIq0m0oenmt5XPFIllJe/mFN/bVrW6dgmflpSIYRa/JzzSaRMp2vrEvY
xgbjaisYyU+kqcNNwyD7p73dau/sbESYSOv+Lh0P+dLs4yCUPcQrwAKNnhMy5dX9+MJ24wT7C9Tw
3CI47XHdVusj5FGZs0+ShJCFHS+ugJfo5o7nEiXMJnsRonXp9VPvPD4Gm8ZApPrORPeAWby8utq6
0aZAJ/emnjXfflHxPkPSrUwUornJEdz0BJ/xL3oxkZ7a7m92AC/w8l0/ueaejAlAAX/aCEBmKXsC
YYvTudqn571eyEWhIdVdpzepJ4xq+nNwogM2uCVFZ4oMlUlPiOtN8EgTgMpbnVpZFdDPMeIiZ9eK
SC2LoJ+WH7VryvHtByJtks4e5iUHOxftMY/8ejtbh4j6xngYo7IDK6HyDw0GjR7JPmcd0u1PcHJ9
CTwsAouSXlh9J4MsQbN6Rtz3XhWCBRGrNDKEM8vlkYZMScwuo2UNbX9R1b2DXDsZAK2lzX/nkIjW
dz08d6kh7gmhOwy9LyZz1ZTEZDlxqJH9nxzQUW64UMovXdxiuP5u0kHePO2PD27RPjGxevFN+tJp
HN/2rH+nSI0ceazKzdA71INoAjTBlYfPephqZP72xROP/sQ8Ima9PK5zzaySm2JreV6aRUZS/39K
4Uh1TGEIVUJ0h/kRdmgCLv5WN4bKXQGNLhn3qoiFqawRYxuyn/WVrm5LSK8GRbyMNHQENnjbi5Jo
TlV/KIupv67LdJeD/Ux4JpLq4k1qQBNI/i/4miqZNaCguzS7l72UIDGCEXbDRO7P06KjwonIAstO
MWlCcRQTiAi6GV/Nqepm1srbLzxAw1DoXnzzsVCJRWq/HWLrimGTQ+O745gOt9P7lp7TMmr7USyB
i7ai79IdNZTHMvUuGTmDtr/xOpgijFj0Nzr4aFzWs60ogLWksjBJNnLVGLwXxLZwZ6E38j6hOODy
bqOlz0S8Ra0PP0Qg86L4hMCJ5wyLo3qUMYR0FaL39hXCv0+KKqkWusZ0XHbPVi3dKqJP9jwvFtQD
HaWVbSmR2ImxlY9DGJ1tTT/I++CnNbMni2bzC4QqHe9NbsoB0kQ7/OsCNvGwzHSz2GzLWAe4MSkQ
cwhu4AZlDZynTgfLAmnfM+JkN10o6Xr73jDVzpydtneIKrq8pNXNQj+p7Sfbc8pyZPHhlETKPE4f
2SZoNtYk0UAEVPrZbZnGtYBEilEREgJYpCWz1WVy3EM+xB58uIikb+Q48sY0V5aalpSmueFQvxo1
cjjmYp84rs6TNthITsNj+EogICdbqLyR2zzHZ6hoD72hthc54Ga/H5dv2PBjlV0TtTqnVFppQmK6
kckX4CoKqLfvzY2k/yZ8kzN9efsngpiv/ciL6a1I90eUFqkr7VHjFESrkyuQOQ7g4edqiulcbdYQ
Z2P8CATwp8Z83c/zILD/ASLeQ91gIwWHpZ0DdleiyehNl0rpNBwMQ+CD356t6giqB1K0CNBX/7fl
tI7vMA0gRl6NKkpt3bOgp9QPU8uKWQz1ZY7xfbrcw1mJq56soes5/c8i47BwdimrE+FJsInODIsn
1hyg+d2gvwe/jArRt+aNA9qTRx0xQnF0P66p+Wrex9FMzygn0V12mrL1tBJ4pNikXXiiJTFhjwVg
0kPNiXy9I+dlB29wQ4jirZ/YG0z/u/d8sMDBxiCyBN2lS4feOUdkG0QA2CR/wwNHWmveVY8skGwB
bEJwRLvjLoms4D2sOUiC4iHzTSGb+5cIR7xdIPQbxV1AXPDAW9dty6mLRFK9iJCe83nkXv/dAeUE
p/A0YWCFLIYJEpIDqbl42+HfJVBLCpQRRfk7CWGipJBjivZhzV1EAh8bn7KibqaKZr1kcd92gLjd
8W2JTtnXUNlpCZ6zgbi7s7NE0QlKa7UGLWN5oL0P5ZZFJc9EAw4ZN+01puEXKDpi9UWVVRP391UU
5xaQJfMYXdd4JxOka8Gf4mCTuZuKsp3HZ/Db7fZhEKwyyGAhDjbL6mNB0ghOGJHTMLwl+o+fwc9N
FmSCF041/oOT3QZyeRc/YzqfqyvrtBVCwfp2KPO2pnP3Li8WKSTefDKNGjE8pS3HqDuQ04kiA3xK
L8Rpd0Zi/HlMzy+3YcgojWguOKuibcdkmIqNKq2WRbVPvzyxyU51mnHoaVs231QEvtwuipY7qjkP
+2WkD5I3VajLFU2RWygGoy2bT0PCbMOc1udjQof1iQXQHozddKjy0lk4K4Phyh5TJLIujW8oCgur
wrGcSdbFaCzDOqjpfAXftiz1u+PDTBSCpfemElmSO8BUeTKyedMv8wxYv/b+ipbxJorlTt66jL9y
2/OnSbuG3IFd2KPTyiax6RwLTE0nXkrZng54khl7kfBulD8aiGJusWry7q+k5ia33jHyIrFFXvJq
F5jf09NHDLbt/6y8mTEPNgukP7qd0/tJKB1zmR6FMcPq1ZWlSe/xq1LzjjmLxCpizMFvqERTTSdK
slLWwJx8oTmYWqJ2JynSHLs9If61vT9RgV/1ImxT7pIdfDvzrmUB58D/BO5JfOxKgZZu3xl7y4UX
kr8R3hLVs/uwBruH5QHnL3iC5bzdJ4q9NgMBVhD4JizAvSU85kw2U56CZZfNIcQBxcHd/Y05CNPa
ITuwIli7NbwKpKy5brl5W+jg3AOpSGwo2+Wio+Qn9OnCNGu/ZKslxqH0PGKlTKZf4yJ8rkJXG4Dy
iwR+fuhmukkvaf8Bp67ugeUVyLQUkHiFiraYAhkZGV4s6cng8MY47igCFuaitTx0ldC3MOot8UI1
DJuA1NHmmtqAkIqjdVOKepp0jPp4G64nN8ZM3wsRfYg5XgZiTn4Bs9rOlo8IDruTlgYduzUDcfOz
b2mDoPVk3q/8hUmwGU39QVwlC2n0tBkgXu0zXlFOft2b6/q8SZ1ALe4Q8u4z1UkeuzNzbZ8hNiac
HJixo7Z9xGiiaRGlo2oCAcUhtuYcVjnnDn8T+BH2WdCS3NcQuRlcmMY2NeF5FZ+ES73DwjhO3LvK
9T7MZaeEaLuh0KHEEmPbSA3rImEVzk+xwkVSjsL4H4l9k1kr0zwj0oiKjtNfE/7/Txx7WWXUHN5H
RMUdLNNyCqsUoIe9lhS4MwQAZ9xx2nDtAc2bBcKJ/LgFARLDbgTItpNj3dm61EfznMXJvo49PuY7
Wvtb+jflJdZuukACqXzPuK8lTy+wApwrxxwx3HJEdOBX+5jekIV+Ww0E5oA8oaF2otGIeemrmQrm
9PE77ymkMrNbOYSkGmXKCU6Ry+L/IBtO+rgWU5vI1boM1+zTfn/R7VMa92sPFtGqI8L0AaMdcb1Z
oPReNQ+slnsIyFyjwPv2LHgnRYY2YZ2v/nrmJcaV0VBmC4NlnxIAN7o0IUhHAeqUXM8JHT5Z+9jA
fY3dKMyRjGdOY0PkxW4YoQbuwIyGN1Vs52xbPmPRU2xPoAPnioDryD++NzNDfw6ceX+10+QJqmFd
+5DI8P0ot+PTBjpdWAvh+VLf2G9pfmAHzDAz3sil1zYO+2aiK0mE1y5zPBsq3VBrvdx4bIwoHGH7
myyAWHMYyV0nVyI61uVyaZyon3JeW5zgXZVW4fxngdn88QSWQT/kQ0YY0K0mbvmm9CeUYl1gHs+b
x/uUw/wxiiwU1nx0ZGF4b/S5IxtQ3en12CkefjUE2k5wipoUiKUc3CrRSYkxNIsTvaHMzRPFzihn
3sI8OmoWeSwXEhzDWZ+KSmDcHcH8CmARHvpVFuc3Y3LRxVevUDt7NQrTjkvgBBgDUio2gM095mBH
tcxg6lRichrr+OhSXVLlh1xI6QqCM02hCDS5PtespwFgjsH7LyYHbmIRKn3+DTDsh5dxp211krr7
oJ6W2LdUAk4iwN3AKK6vVpUbkBIXPEHdhCz4lRbcs1M8Byjd6mFeUbZQrxYm5hLH9HgYgXLZqjj7
eBqCjla9w3CW6NPTjU539OdeZS3jC1PDuf+cz77nISNddWdX/3xfCoW5DhD4rcrCOROZ06efWYew
BFO/5dhV2LaMeMyB7QwEAopIvPHhU8HjC9GIxUGm1zsp534zbJCFm//YQHKZvaAc+CUdNJOACATd
eeaet0PKLe+v8n4VHwzlsKCHj4QUXlm2mW7do9VZ+khzfTGJSAwkjHUrjNxGmdB93Un1WLMTWfN/
9Vox602/N6cuYQ70W44HGPA0AuEJQkEi8fdEvKAlp8cZmnlkJOiK3GuXYTcDMQ5ikg/HdnAK/dq7
IEZvDpz5fapNNyCEco/v/utLpMTEoBb+2tIz9MQ9aBDLquItTNjd6Acvamdy2vCi6jFC/PcxkoHk
0MIGgDsZ68eSww7Is0MZCr4mwEKBsQ5WaSL1Xq/DeEzMjJ78Cbg01r/ZTax5h0XfOuxbg0bnMgas
g88TUgUXRqdd4+wARJSrfAjvSNb3fFro0aq4LRY26noB8f+MmAIhQMYl9ytAOs//jfm5sp/meOSr
mvTtfpWk7w9eIYqJTpByIy4bpeTuYtpLFQsPs6r7WAaqPbekm/J7M8KiTHvWTv8b+YhRw4yKt1R+
G0fh4qdUQHor+cEybR2lqr0VtkjSIgKwuhbExBwQlq1JFgdpEpWPo+SDGni933yD4uuGrJU/h6+g
ZDUZtqcq+YlLa4qoGh3+If+TgW9CaE3Na1p+WUj2eSq4C+KU7aOHrWkwqLpZqIAsB1M+RXN33upp
2uazZ/LXlcmcqfcomb9hpfir4WM/WZ7nvBnUZcofTa/QkbWfJW3OFiyPWsPx8CtpPYVsfdCkYSdu
RZfE5/q35wMjGvdDX6YTJ88oc3wLFxbKCh1k8Q82kq6wqMiSgQdADX2IjLurdcyGDPvf7h/Nq0ZQ
mM84sY/uPfQO5OiuW8YlxaMi6vQG0iuyOrdX86+T3Ps8BYlwjcaJeAPb02PlC6H4qrgy6fy2fZxP
0WyeVBjl8B/4dGz3xOcPvkyTHu3IczhdqJBkmrIABHXRohjkhDa5fnmnmGgfgjISZQKmCg7Ub7Z9
jHtDqGsNzM1inw56FcEQQytqmkIkSxT7MOhRZW8GuwcuNlfAzOTb5dQYvSHunWx1UhvhQ/73/7+k
FMrFqfu62DwvnSW9HUTb4jJya0AowEoiEQEN+MNdUODO3kXuzg3iZr4x7/gMmf5FsBoW4bXXHaNo
e5KSHPQqWbrlfu4pfb9St6kCaxbxDKI4gpEc1njopKJRlpvP1ktUlDHfEucXag7+S7qD7bq4fTOU
ukf4/Ck1NlNW0AJlZp3l+3JPozT9NerjBseU5+Csk8j930s4dbpuB4E6agfnA/rjB0OeojV0y9Lz
LEDUJvforso50fZL/SeO78RTISIDjc1l3Xcg+dqYtRPQMapQhddhqC1en07B0i3Pc5yHT0OOzKKP
5FBrclssIxWiusexyrjVo0N/kC1SZl7jKcivAB9iSGqQMZfVJg7nTMAVslS1bN5DAjaait4ghOUl
5SYqjvqnk86EL0F8Tuk1RB0MPYRpBymS9U1U3Kjf7PuwNM+AS3ilY3cZCXuB8cUFbAP9+2bcuLUN
Shl8davYLwx3mBOjZFlgE5s7tFurroRGqgRBhMzmo8du4Cfq6/uOCPQJny7Ly6PYo3r+4wmsLHkk
UBgtm7vU6nhqIqya8t0i2k6b6YxTBPKdf62HMkInhKySv1mIzzEHxT+EVCnxrwQOPHd7JQ8upu6i
DMeBK3X0D+dEFqOzIuZkp/6Naki/CM9r3UjGgXEveRExObvEuvZgp0UK9+zZPwI0geQhFYXD4i/y
EoW1D/tZrBphZ4/8J1ao1Rnv1IW7qSLirNoSvUKhjvGY/OIS/cEZL0CEHE/jp3igcFCXScxs54qj
refumX2Ivbz7PbKDXzAEdWhDGNXrhuvjosvHW5Toiyl4nKFsol9FnN5rJ85Ca3VFChA1jfvys6MT
AYJtxdbseLCcDRXfBzuJQJl2u9tkHdhlpGJu3XzQSpFqJzVBYrReGdEeBW/vbxacRHQCtdAU80x5
MYuQITZo8YhDt5WMnvA3EzmHS9riLtSQaSFfTBo2Ar4tIIr6RxcQgi2iI1h2EcNHNrOb0hTtsJWO
O/eah4XnREZc7/z5aE5AYJnJ2nBR6bnS0QIxoKraSAa+qMZ/0LWIQPqGy2zaUrSMeIcedhGzHXrl
R3QszjrCzuxgabwwKRSP4qPPRaNQFUQkSpLL7+aC7PwIOyFAWe4fTpqmFPtXs3xOBaDpFnOA3RwO
f0w8zmBFZG5Q16ZOCovWr4KJm6kFMSLACN4o2xOPZ5rGKkEzoTLDf+OxtYhI7dnM8N++HP8ADUj8
c2lNwhAnDqu7PMJ6nUDt0JWtBNdUFWeP3QgHBNdVfzT+5o+gl4uITKnzNG2970UKD82v1hPenTew
dIgjnFq/YxPAVC8h4OAEngQbl1hQ0kZo70Ouod/13KYrhlJy5IBfadtOgp6E1XcCmz7OwETe/F8Q
NPxcLt+1gEEbSX7sGOJLj0JvW5hJ347CyOA0mRUUEaIfXbFQyIGCUkidrX6AdSZ0U667m/ZnnKP/
la11TqYoJtOi7vtZmFRLjaoH02hRU/xu8JmR5henvsnAJoNa5OnPE301EgADyip4yQqGYWcX3CQD
6knzHS/vs31wa+SLj8/ZSEr1v8epzcSZ60ZgrNP1K+ttRxyHD8tsQbF+slobEonzAxAfJYk9QrN/
GPuPilyj07Urg4wYZlGx8ZxgXqNn9RlyWUhLrEHAIUpeTGYUv82WaIb4Fzz0leUgu04E0CnYRk5k
AmJ/WLeBA2EsB7dB+XaHZcNN+2LxXwHLgJTL7sv4OkJZUDNJACBtDbMzzwNBxdGwoA+a8fw2eyru
fEAh3pt53zp1ZcI1HzcsT7vTOf0Pi9rbQoDxJd0/m7JahrwPhm8fR61HOm9xBSJMLGqmN3QX+13F
uz2nLY5TfyNZ3lHJV+LdVXWRQzzAr01J4WW8I4p54VWUto0Hqkdv02kG0jQtR0jfebIQgPFXbO7Q
ZK9gNiueRv1/DrOg9frxA7F7C3jJQoODx0g4A8bRrD0yGjuZGWXyFChxZDRMIW5XstF4Ogh09Fc+
m2qowXn2slH9zoZjS3dFqm1nDBFrB3jnePVLgmRz+O+EXRyjo6GsP36jUR0uGdSilpTPR/siO2CJ
GIbcbk5yUFG1ZFahP8EfPU+jEt0jqRwkSsLf4PxjJdwrFa+ahlEN2KJ9whj41YLse1vfP9bLAbkz
oYh2ZrcAVPlthpj2y6EqccxRfVsZ8KAd9jx31Q8Zr+BkSB7jPyIyoK5/4MpJTpYytn4/klVqOiBM
pe57hIrcpF4M5db4QRpcWjff7atMC9zLGHwdEqqq8QRbdsLFeRQelx935tJZuxOXQH4hZwGRmnl1
p6cook8gsDMiemyXOYhO2ohv0DBYSRvte0BZLkiXCkPKc+axGdTRnfNxIiAs5xUPIpWmREJ9HBX/
x4MC2L+VxwQcO3iQUiOAAbXSWEYvsm8FkKzDJp/uDCue6rTQOur2iDj+rvKMaJGWEQLIKp6CLFL1
9qClXNdzTl7ZR6ply/+Be0onB9DCK16yGBPFnzvtFnV1P/MIQ1Ld2mA7HyWvom7CfCjr2jmm3/sC
aPu7xoTJvLBt+GVgJ5Ez1bG0IVbcDKJELXsqPh5DGpEx9Pzs20Ra/m7qaSBh6j8SX20wKHOazVY3
sIjAGeaCy9iYs5qxYXQEnvvOfkh8HUsYs4GQpJHeZ2fhvN7WHLBvK7nMNeLizuy30JoJ+D4ajpEK
PgDzfM1l17r/x/AosNduPH0/cZy6/k1Z0B3H6ZcrBRje89yVCqPo/wb8ojQWYx4JW5U4DEdfsNHw
9RNWBjMw/Y140C4APi2NvoXNjC4Ec1lrMsX8fDUER5Hpyt1o1NKIZjGGC1qfBs4+wCI9tZFCI5MP
PkPqWgGR2oPuo1frSOiZE/iGU1yMwLSTZ9zg4/a7kdRCJ2mnm3zldmk6PK111GMe2tiVinlf1rxm
v/A6WEvyz9hmirkoWjZdmocNxcLnk2FvwuTeuqgPpwB2NJCFAol0/0kJrB8mCIhRyYEpy3czDbCQ
W9bxGFccJD9dI9ZcaUbWlf9uqziQGZs06FDyOrwodKJUPYAAlzppTmq7P49zoH8xq+B5HoOdOiyF
bqNYcAGYp76EpOEhsJGJF7MGnSCqw1e2/U2DMpfcTii0YJNmwuUjw7svZMlbvj7SJRMz3gUeD5AK
Or+i4XUTzt/fLLxF6N00jehvXuMC7mVdJzX+uVZl4n2F7N1KXIZ0KHXnaRSLA84uqtP5dem+a8N1
+rEMBasypFUJtMPzHwBltA74qV2YpwTA640hoslUWRRtppDVCMmnYU2kBsXX/nclT4wKQSbUxLDa
LZAYNIII+8Zj1cv54eu3kfDhkd75k24CKvs3aA/ClbBEr/gAAr2sRePeby4VcfirKV0vLBesdBm9
PMudFbWXmYmNh0llZnxfWLYz2h8YyUCzi8YoP9+am8zAfDOSLESAYgmjm0XtefLkJhGmL5jZNkDb
tIIdw2we4y2z7AkORYn7Td0ORsSL20PwnXkKVJgW5JCDwqG+CshfPYg2/ZNRRmlPUecllYCsls5A
k5VFP2OPVw4KQxevfmctVCwGwWfi3j7s1Ffn0nI/4AnA6aTBRS00ol2MPAsTuXWvNAoiRabXU7ao
HbemwMsxaete2E8iV4KT9QBaLoeHmhhNvEhH96cUVxsExOPipuIZu9hOpCq/DBq0cwHZMAqQTTJr
96RgkyZJMZ47IRwHGbXVtwnsF/+3hbcEQ3mPxrKtlc4F7E3cUqKXEJnyA3iBPYKnqaMwqkV7QDoC
yc6xB0Z3bUvSBqxWhUQ2uAQ74GVIGvxh52hc4X36zyhl3bQtQbj2bWp4+tQBXeOBELMk65c7C2lQ
IFhl97e2gwhGcJAcM9KyybckWA/A1Vt9ABvR+6YEYxZ8rQEhzL9z4zHQKcvN7QxSouiFaglwf5OJ
bteLerxMMfk9cOjSRAPP5mQtgpP3//4U/PvZA+W4bH/GaibKjYoaPAzo/lzFd3E6tr4wG8/mPak0
uzxEluoKULq8FEkuqTAckzr0RnlgtRTJjGrhu/NjC2CBcGb3OldUNxCvyopi8zH+jJMMtaqUrHAm
P+Fwa5n7kFHuaQj3FSws1WM2fTj41QdCoeAu5RBkhwXHklNYpah2h7tJDuK3bGUBoTa9yzvHWska
7M+GK/XEJmH4bOnBeEWjnPZnG+6mrMKLT1YbAlREVpcjRnkQhRo+2pjdCl4UwjliuYi5b3j1x13E
TlEW+BqY2burKXzx3iDY0ViD9cQ0EPBdHyqSX0QWxI/r3s8+42lmMFvLLFblbFU21ixkY94JjHDM
RMcS63+d6mFtXsFsqRvfNRW00Nx1Noxs/f+os4gK0iJBE0pcDsqeqq3e41K5XvS/1bp3RR3GiYzI
TAxI0dSqJ5v+Cx5CaxX5M1EKysk73icLeerab056BOVpJgSe4u4KQF47xbJzOVtOSXY1tqkC3gxA
OoUGIQfqThRM8oRp3QPV7ZPOgYp3setchL0UH01NHO0bnFT/JYWr7M30Owc7QMP4V6EgxOZdmk9v
s9PjRdSdJnznXQeBvE2fwjkI76EoaseKb7BQ+1TPaPyGHsBxAsDgNWA3cg4qeUC/U5pkf2ispCHj
dwm4/D4oJISdesJoS8xCkerd5QLIc9fujCG7latfoW4cc+7HSbIwy1CZ9H4k6co1Q/mxWAi1Wc1N
tNYGT7UCnFULJc4Zd/IPcKIC1xsfgpEnlVRVJuXHjJoZMo40EbEwE5EYNKcT84HNohFyQ46ZNnek
gaAaM4uN98HAD8GDhC9U0g/P553SLoHu8ald3o7L4c1xCZiAUy1owKIYgdLUmB8W1TJ7kkUWA9ej
TgyVD7H5BgWlmpRBGcAfWcepMhc5fSvdmhll8NoSwKC5jmqJ37kEXUXKTyOGBzowb578L2K5DJe5
LAzEgup0FKiZJGD6NmQTapzT4tY1xNGUD8kWMvQJWbCyYudzjCPQJmLMW0a2pxStwAYtH+QxbCcW
85clHnL1tjs2b39QFBr1PJrBHtx4UaJlTB6gkxhbQFhm6p4/pc99KBYR93Vbb4DSNOwUoupA8IUT
ECvZm6mA+Fuzs1/pd9lmc0RR82CY53N/vwiVBpv7LzVIKl+GwFY52f/xyAFpTObyQwjxlkcsnC/Y
EgxEJbEiuxGFyQvE37Aqb+3llr6wXplZ5U4CNuXE8rIBnv270no2pRDjoSCIWhGTy9onnGw91U7t
oSkkT8GS+eljHaV/rg7Kzyh/7zZuEs1pOeIcVtsOexeIYjqr2ha6PQ7iW++ntZhe2mhSERkoCYey
+dbmS57FKpwgua2nsrb9isFlI2D69uo/vMml0BvpK3J023DeSUwOVzOgoXsj7E7/DozYZRXuAUSy
bltgDjOupM6qlZ7fnCpKzUDxzej23MaQfGeIs+lRtU+XPl2jqeub8gVcGItNXx8hV2A80l6lhhDf
dj49XIXns5u+xX4czapVnm4RvVYLIESPRTdVyoWNav1U99mwGqandRjviChTV1ztNaP1pabqspMf
g6c5CN7UoiujfnRPCHcp2Yc+dcGC09EQuWQCYSOzg6zeIwtbtiQbAKnFd8WV/oWK+TrVjRFWeTaw
oKbyCdi78YqhQOl7iQDVWEZqrFxI3mbkpsFw9o2PX4bb8aiSwmpGi0eKA17xGkuxzm3LIUxa90qU
Hf0Azy1VqjiGlswjzhSyJjsWPBVLO4c57iYO4cpxxhNuBAudpDiE2x52l9iGKZLi2Zq3nbkfg2WN
tHtkGAATbG7fw5nbtLZlPFw/DpBfzSxKp8rQFNDjg5+IsFpYNb8khxVVrTf34UIGndsWwJn6t+1N
JEnBDxzYVhidkAcNEU6PkRNXnBHsgfGL6p/Wv8zAoxMUueWNb9FAwBfQ+0fs7OY4FK8tvSaF5Cda
m43MzcBiFVTlRRLkpW3LwkXhWDsDjXInXk+77BU0IX668pd41T+8+qL5nAeE8ohVbYCQ/8RwuiEe
mEeob+6PZ+Ti2bDv6UIXOyjvM0tIa6WCWsGeWSDf5XYfeRBzBWqehiGPQFOzcFtExVPZKbfZgjWT
EFntZNb4JkQqpF7PxpPI8P2LzIVv+K1eoom8mH/jUvnkXemhaPhd1ZyQ3mVUnmL4MVlDwHpxZWaZ
caMpWTsjnoce2endJWr7im6suqLTpcz91RdB6hpN/DzVhockh/6A4Rm0SUp3p36ty8zgiHgYZGel
GiosBw8lRbmAnN1M7+i2Cc86uNX8+P3A6ZRbH6X1cHJoUcaOPWIqVrBUTTuFUcquDxuX6Kz7AcCt
kufGI64E5GjhwEmVf2XijTKOITW5dpHovpOP5pkQklpUWqE2B5XJ9vTCRMD3+Mupyb6efXBvuOC9
xRftqdAHyWdyfla7JcdcRB+Cmol6Y8EPEGIIAESCHd2C2RykiLaIyajcSzUNStc/Pn3jc343KJi6
FhldKROEFUooFzlpWFj6l5M/pvieuZfPBsJUWbECRlHxO1jjiRJ+OUCoIl3xbRj10MyuR8DIal8S
PvNEDAO4UcDwILPnHmKex4Vz07o7Cevx6bDQORKDlR359hcfv0l36ru9ert1rkgoSWY/16C4KVfW
Sv+jrK3gURAro2gBwm5u3TNEPI5+fwROStVnF2ERnQjkvg/ervvig+smW1VCaAwTDFFSXQtJcuCp
VIKNppmoNj2zhvg/Ina6EAjruHPCpkCeuMSWp6opt2r1KmWZoksdg1TPtJvPSvfWl1x+6gP0a1ok
XO5kZ2q47ckD2fmuxypmc1cN3HnRVaJtaGsLl2hjxjUrht47Z0qZ6pi0lu0otFxOBMfmkW0VKpci
qyQqjQrz7PNzlRZy38jfGFPIkoIbritSTVVwhHJAsbjPZS+pIG+f1utIVsp/eRwztTUGyBqzjRPs
WhtygCCAUyrSFz+5z1Xa+S02PxEvWac6VCxQSHEqLZRrpM6p3zJpSopjHfQ3/Y82BNzP7ehCqg76
M8unfHWnHYtd6K5tAC+caIBWVUt+9u1hIB4rQYEJhRwQtNgsI+8dotYfH05iBUZPlpB2mOM3vCVP
VGwM+AQ6VIMYQ7HfImsawcUeiv6Ju9d1seNYsriUbmlwLcBBcZiHdw9wEpJT2F8QSyUAHO8ZJpJp
6/+AAeEA0A1Yf8PD87Fddx6pVK3o+YgSX4zHR1MB0DI5gH4egC7xCSBy4BFsZGy1fmulzFwY34Da
GIzA2EfgveB02DMd8jq3udNMX+kKAPYgDT4YZlgMk3waf1JlWTRjpE+WlZFwRG+M7bbHOZMsH3IJ
CHq3NjLnqLtk24kibgKFpJrpi3NRCJeupvfzfq/h9jLGbhAIHvkKAWjnMtUsrCDI9O940RugUzxr
GBugQlnBKhqnEdoGQb9kcCfEjZ/aa9aC5k2gNJM77TtrKwOOcOvcWZed7vcn6fq0ao3kR9DeZxb7
LjrvZRucPRBlq/XFQnw6HM0GHqD4+BqAXC8motdT4V+U4ZTX9cr1VZ17Z0XZt9LhctwoM4rOibUM
X2BzaWmqSoAogM9AEYVeZO8LpKl65wvMJLl6vBZRrtwchRSsqs172V0TNzpIR/iLRuf8zsvenAvh
CjqZxuEGqTwSboGD0Nh2DoimFmf5T4FziT1dYMZ+3ys27bbYx++dRJNpOFcBtT9LpZBMSq3ECDRM
ca75M3VI/QbvGv/K9DqfxcZ/ZSU/6DuF9xD7a2zgPQ1fs6xf/K+3HP45YSHuTbMQyK9eJSJOovMr
ZRzZjbq9+l2MbrTILQsBeiYlZlX058ak6sH8V9N6MBuT50Tq6f7ctuaGkCTvOxs1yqhRhgRHZGaR
5wHgr0fN0xtjO/NEL5qP40kV7fAcjTWMIFeUZBJ586c4f+hY56UjHDfUL05Za7MuTmQwHE+gm/ys
7X6Nj/NTry+2n6OPdP0bVbF8jsxvz/Fa2ISJO19mInYMjqN4UnWbiegDvGt/mg4QisU5W9QHjaJ9
WxK876ReZ7Uw7Soj8B6fxMphDeqGTZjIEdLwm4xilb16y91eRr1zbUmSwwY3BcWEEdxYgyM/cob1
b4gOdAFHDpxsCntELoxUAj+l51nzaIgPHOYQlhevTtKRTXPHrSb8iopqZSXgUmzKT4mnAk7HNzpq
J/OHydUAQOHSDJ1nsQ4NQ4D2BLvzB/rhKuLEekEECiCYYzLztZeD8Z+314Nhkn1jVZhShHRyqfme
lO/udREYIeMYLQfKsTIleSedKrq+TfwmPTgNocWSiDjc65pIKwAAsNsuXvJDoMrgdXn4lBQJAZ3O
gOJEK1xDFo/p16BcHDJD05sJwO6besgPs3ccjFHibjQ3yuti9LeiTPtgwHvHu+gaB1Hd/9Ryb1ll
mRfvTasfkoJNXyGDm7vgXsv+EIVvHRoC0yJ6KRb55dkethaJLe1+kBytFdVXoT2rtlyEOzqkHjXU
KaWOF/ZN1A/t3SxcbYReZS5hIEafCfyOqFUOVJijNSgEmFDnvTLVHZNnGuiTjR7YBi6BDrasE1RF
tW7Yhgu1Q5FznPDtH42qDhe+Pgk3CvCHxYRfwcUhRJDHeFAmgWwOMK9dX8wv996JDspdwaxDyfHi
42mSFYpnT1B/NyM7y17bqCobjnXtHTcNRtaTy2YAOg8jSFDqKfeNhoGjBzXfMsuhyDEvLyXYJveh
zsnll7VrsKepGVl8ioC/15++9RWTomCG4Ne9yp84YNleMYAx0KT5NUXc4KPEVUNkVdLJlI9iortc
0wi57m/QrNFDBGgmu7B0ZKbK0lik7c86Q3VlFsESzey/jKo4tnfLkVK02LgEFqYoZsaFDPrFzDiJ
0IQsh33yJUjS2KWJH0QQkPVulXW5QS5XrdxFlPunElyeZoWlvm1GZV1ePK8TZ6tj6JxgsJH6qkVu
qo56kZ1v8wcGZe/sV136fwrvif2dgKfxBk037P7mOgLNRwneB1ypOBpz1LBvS3APDORi/AArs98l
m0TlDwl/nVhIY9uvo4fxuoKhBe2GSfFnCyb9vhFhhVt58GvNlty5CGSmO8OVNnUb+trzTHykeEq6
eC/ulgBo8m1zv4LTJIqbU0JHWBpmX5iKMThwyu19RpoOoguhpiUF2xW+7N3VRotScWb6Z1WA8Xte
md0BYCQUksGrxd92JUDIDxO3eEL6hU7gtyN6IPl5pBis7h8Ya2gjgX1R2+ca0ySChUJbw/psfIQj
vR14Nt8xyttNrcp9ShcXfVkufnp4uKmhG0gZK8Pvvhkvj+vlYWXw7VIWNiM0PWroZ+2xdg9TUQMJ
g2KPutBCOn1ZxTWvp9z5lDRV+o82khfFMomjCYeKU9dnV8sm6Lwx0ysArr5Ff2Nt7BvAaJHZgDFa
YLHeo7uOFN6x5uC0kG/tr/Adx1XNj5Jwx+eOCOpznxnJXxJqB3UIuVN3qLjIB8o7YGHY0YQa+Zn/
bDn3eV/TqrauPWSR7sfrFvLXAz2dDO163Hj7G1kzJRkznklZ5d3sYZFqCvON93dErM4eXPh94Sol
H/9lsqPeyr/cgw0zvcF9gmdn8qxOU1uRkCVQePB7wjxLekmqjyoJciAkrC7pNVtgFG7dYzokuIL3
m+prsiS540f4MJuNs/5lZyQ0006ubBc+MAugFhRwbVNXtusJIa4CensAia616HNQqoB0YI6NYhML
IccJfu7tJO4NeCrAHlZf4aHH4sQTf7KPcReZ4oaS20uwu0zFo2Z0FAkbU0BgZQBLFcihusfNUbqu
JTDUW9et1rwZqQLQXClQ7U1wyEvI3F08WwIc+o29ml3+48AIVDGKoDkVhqLrjbYfOk5YmNp5yUB3
DvIedpeyZV2+irt9BR5wT0huRecwD6ZFuYNw3JzC9OUWLu4A+yMCli21YtY5KY/SjYtSJwYzgt0B
VJJSCBk6xSFgB8ju87HH+c3ymIcuZss/3g4aVZZ39iOiZ9WmowOxXEDEN/fRryJcj/F6vC4ANb2B
gCmLPFtz9vOXvDoYU+i+UyPs86psrhG8P9cVfVeomOrI0VpdJQLNote5UAfakwu8Trb7jmV/FtyT
n5Quq9vjlGQDS/8XA7Yprd2Y8uuA2kXunKvwWT+c2qJ4N3aRrGWBABDUNxLB4JP0qOHOxX+/48fE
S0FDnuo5BnjA6XGdEjIwc841IA1MDQOuhLY3iIDR2j1Q5UIloU8+KgMzDu0XXKkSqs7EBP4f5509
j83Oaea0IyjQrJ/6hKILHYQjMaCZ7gQqQG6cW+NFRI8STvdXw28Omdr0OTUlGScg8b7VypTIu2l3
emfPk5UV7WBXDWpQAebh7FqH+C3/3YE+S3z7ZTd9XFnF7rBv3OzDJUu7xFmUCzwTHuOgl6mKTu6q
qVN+E31qkhwG6rpNdWfASd9CeHaWmpi+njnUXMmym/6mqsx4vuMDYMkzvuImkb8RamvOlMeOTkbB
gzs4R+pqWn+5miNklpm1PXE44GLvyuRo6K0UqpAj1oioVNzn49jP1dW6I1/XOa2C3zzy/lPFOMYw
KGcWvtmvSzEeHQFvxGTibiTnsOYk+Fl6d2tEQzDo+AS1qFZ46JrVSRkN/T+q+TlrtSVwPg4YrNF+
lTfmFtcpapIdEQ1XcTO7dmLxIjJJK6B5Unh8vexMwl3FdwBnskH46PTwxWttEPfMuvjglS5nE8XK
xWy4oyORtyLOftUD72qOWHnmBPUGml47STlM4b55P3kplLu79Gz5tzZDj2UDHfiNvCr96k2UApHv
SR+SsTsQmJL7gswfKze3mI5edXccSlwUf6f6e8+OD3PyMSe0zTgrApO1cNxLPL2bKeNUgra/3Brs
i328BRZm7ZqhOecCq9eqpkF7DPiIPXEgkqfmnWHixHVUEMzaO+7wVyKd2F6JD66bc3PMhaNPEzSo
e16eGAJUs9C/n9qvBe3d8WHuErI8mD9EqgVyJg34TxESkohk2BYv0fhHOf8J1cHE9JlEUJaOlcqt
3W7FeDOseWT5DFCT4ZSpRa7/BNGggXaGE6wnvzmSBVmATtNULmsTuyFdVggt/hSfG5iCDLgv/oiY
koF7fTpbqK6i/7xM4Cvpk9iZfvSZb+GQpjY3lHA0S4GSssiRSGB6wq8S2hgewF32fbwBrWr67wVm
/pqqWX7imv6h/5Do38ZeqCbNLD1fB2E/ySgJC0c8POLwB9zPkvHMU/AEB8m2LjNH2VkqgeL9ssx9
Algu/J4Z49aa4xNrj7o5SxLP6f3SK+X95WaR6cyRnCNmPw/ohcZ7fJpibcGzJ2Kr79/gAaCbCHfX
hZwOUx9GkEKBRhJxrJEWhsn6L7+AbJrIZ+7sXpFNW6rLBOin5wHmXLru6kcOG4GAKN+O4JUS0bAp
GqIp9hvn3CIY8UcAEX8NB4xucBWsF/qBNbujHEaiIndWbJ60y6GeKrytnjGME+QDpUtnSnkb0GEW
edXfaJTAU0dfaLttOK6sRg48GEzrlGZJkb70uKaCFWagtXXgtGtZivv9xy9GFaa3FAbTqNUbNSwD
WK9uXHDwoRasJp0fE29OUKgLAvzOQkzXcAtZ7+ftRzwm3gpFKbvspy9sTWKtXgyMHPOMt3HlAY/Z
4nWtiWA5STrOnqWpA+ZBKu7yem7I3oBi5Fm7mK3v4rqjeSNIeGMgyJjXHgMcC3dl1wlO5PFodwh5
P8rRywWHdeupHNu5g0USi0FxX3GmKthy4K52OMtassztg6Si3O4qOP1zUW4jR6quF3voDcjyAMfs
WQtOlIh5wsEsPJAOg9NkCl/mCJ1LjSsxIG2ct7LiuHVXNOb8AQPCj6HYZKCCYSYawtoOC9utpoH7
VgoudGEuLpwp9mxhEz0bX0uf73QfexzFTMjHEKE3Re9/cPKhCFex7+xS5lG/1DA+3rDSk5oYUfXX
oj35OV6BGg6GsCL5h7LfoiFV9xA0/RPdz6Oizd8Rhf9qUd9NsstnSRqvvOxHR5eid6c2/g3Xu0Wj
oyEH5NMw3poeXRJZk8AYWfD2g431ri9iGpwOIb/UVrq4QkON1dNBL3k2l/qmzhVzmy0TD6mh95MW
XLZo10CHQxvbIqNY6Q+l+NEFER/oTFsbo/eTFKovPXFWCmLuF96VNGJ5huNUZpUaJPAmxI3a6Hxr
6M2hCRrcogf1E4zG799C4nrgT6b4PaQelqGbE9H0XRTVr/M18iSIfA4V/sxLr/y9x5Zib4rDPsnv
CvzO3ttnyoHq1jCyxoPGNAqL4c3E18dlkNSLrYwYzfWoosm3T1USi8rcG8nSUEpNyFnrWCkjsy2h
XU8kuKgpDjZoS6Wjc6x9guhrJSOlUo+s5capGlhOGHx98nNs8w9vpq0BZ8hAeaoiw4AlzG1x65PW
Lvxm3xNX04TGYfmJ/UBwi4E1xaLKTkl5SF6DAKG0LyFI88xhfpcpDs4SKBeXT7ZJTNrUqvYZ6Q3P
GeonFUc3XJ6WivCBob79e2NSk4LqCq/kwpfaraRS9ozoQDWjewSyKuJp3rah1nw4fV+0chP0kuiD
FDx4jXK/e9LP9u+S4JkZfeTOVLgn2JvMzTBuU5DOAcFVizV9sbzBDpIPtZu/1i8a+/qoXfzzM5/u
IaevYOHFFT5dnxzoGsZGdmUvHikIASZ/RBL+o7Ret95kYX9AwXN89qVbegfc3IZzcRv7htcCGgvQ
ILODSVDL+rHAsnMlxjiM+8IJOv32Wz8Br2iGlcXEjo3rMYfYPZ3HBCaoDZyqP1zOMtJIRid8D+TY
yeYEeg0gh/Zc+I3nA6ZmiPF/mWQUjt0bLZR+8VqaO/uBARvHVSjmwITLhOSPH+T3i+JV3A8bgvX6
tPIhzy8yGI88CkTxlUSr5yqpRmef697brodo2BPyjuheZQY2Wsz9lrU95jji01CMZgtVEdaSEqME
24WiMwaDTYbB9DFW1iMdCT74V0N5K1gk++etWt++/0kqHBLvd89QvE1vzBtXVSFG2QE4lUCFtSJT
rUXlT1IvA1yR3qW7gI3cGvHzYeiKpH1VopJFhmWaISUPInzfpbodmYsD0pLWLCbfgVKvK1/g+xos
ERWWuZx1Jt0YGrZKeSxt8aTptZuehSfo69mVy3yy9qhDigwy2vLtURnDXLBpf1e8QooAfh4Z2BrE
+Y7WgItZnK7vo9cpzHUKuJjDCLo+U2fgtMSLfws13tjKTX2kjDPyCJ3a/4FGQXoIm63bZ9msFIjy
eOJf18haFwv56q7acwLCe5etYjFkouyn8i9x7Ive3Oti1PyFw6DhJoOphHWfdS7FV2nwIf6qkVM7
U0leH7EKzcqr/2LOW0VkNJvb+TU9aezOfrshoXiMcAz5H9lnT8DQnd4kcgctlH6OxTbCRIrdjkDO
yjsJURCbnGDbZSCPMSmBW5z+ENYbO+Yi4sOesWiAbGlnx6Ol+dFJ5FZ7gNQxdkTXPCPROE5PKuvM
0REugCXRn0ldqE67sqhYaTtkNq+4hr3GNydSyDJ/PQKcV4abGi1sKAVk7f6uF076dhFFIteMHA8o
HFpnihQ5CLvT+Pi92rFFv7LRNumZj01kmCnSlhttx5wA77fsVPPY+viAIAazgQf1F7tIEs2LuVIS
Q2JOo2B76Zx+WvW0hmZ0h/+kSqOEfLfFjoIrq3NqTKoMV1NP8Uxc17ni7+sKJJLtCCjz7VfzH0cI
lpe9ziyo3GDafsLU75N9RIrCi4452o3P45sPHlxu1+jchrW7tQ8D4Zo+vNE1xFyhRkVpVDM7sMdU
lptGasTJ+FtSLxLJehqKPl/VWoaR3j7eL5bY4h6WLDL/PXHlv4JDCstdABmDcP9fCgDuneJu6bUr
52u84tqrmQk9Kua/5+hO4pDq5ICQqwZrGQ4EYEEXcI2hAVcosCDt4ng9Ve/1ds5s1zuHaEERtIgy
e32QHDP2rqDogD0pkaGXJd/4i1R9HsFxBAtGGVCe8km9JnkrD+FdD2uC56c1G7XDOFE4Zi3NkbIq
2Dv3W+eb9KvHwXNUjlg1VaFUP/GRS2bBvbFBsBvXEYreOHW/vq5tI/Fj2cABASehfAODhARscGmt
6JndDkWUzxQXhImt7w+ZDIWQcSc+i/o1HpZQ3EcwsgllkiW7xsu2f1dGh332igoR9FkMZV8+Q2py
OXJJBOc+B1I7h8TPxLIaaz74wLOD89thwE5Kd2KgMIgIS5QE0YsVY/I7ziXCHrKfCnM9o1INIobg
UqdQgw6IoHpRbxwqfBSjnSl7/vJcT3RsEKOv39W42rU7hLO26NoggLoW8hiLS7x4cUmBRDYEgg0Q
c0FkTUMj13ksZUMVMSrCf0gMipN6ZkGe9fpOLQmll6HDyG1bndMkqwpHVJn8hSvwKmouJka+iA8F
vWAvpZDPDiEBtoFD7+IFuk27AdgZMfWx5XAFGmbCD9jwjjgoBR4FXjLgNrTL68X8j3SWmNf9jZ0p
m8RRN98lhOvw01IYBXSNsogQOP/HB4yZ4MZYuWwj6acNd39x6KILwhnhLmJbiX0rtjDnTorYlcAg
C1cVYBIDSh5DWPjOw/6r5zE/LBNTEijgbtglf5S6c3aeWh/h9bYDttgrWLA9WBIfXinOSfGAAPCk
Lggy5yG7bqppL6rXijn0moZUoh6NBbzed/jAVHD3x4atOKCNnL16qbWZN+ezyuLHohD9DKwbggME
siqYIGqDIRnJexkU3uAezph/vAdSnpw7JAMnfvL+Xmf8PgWk/MVhKtgCIIu+bSRUdeaDQmTJEVql
E/LcY3lVsUQjdvP+AvJ5Z5lWaZd+YVvgizfo+9tAT75P3aOZHDqDhzd/sq4EMUEzhYksq1mA4DGK
9JFfBK9jPrIrfclaVqtWCQP+ZySEGA+njJM+2zDZBviXeagIrP+TMJbG9iyrZcqMxpEI1t0LHQTb
OTbZTgmqWGWq6RtoR30luLsc4fMcvkC3t1AYBpH3YEhjXFAHMNlq+fZSEXpy/tOIoU++ca62ee3C
+J/re9rnxxbQ4DUTRWE2LrOU0IpP/y9TCYzGMgTyWJK+fU6C5uYfeDFNPmk5dMDDfigA2RN+KB87
Tf7+lzB8xUg1KRv90Ei8Qsty0hmQ1qnIETF+pEpjwyN+lhpKfyXMzg2Jg/CrJNej07mkD0yRdeSV
+/hrwrIatiNmwOv9Bgm1vdzcz3G+2AbvS9SRWPUAEcBVrtGeyTE7UHURs0uJB8GSJEnwwrAzLemP
HrdCTAC0q/m8/SGZLoXP5iRl6FdACzt4fGFfoa6/a75E4TdZcdJgJ19NgwStHUKuW4gZR3M9hR2h
c6zEwoa4mVu8kGucg/T8cqbqMNWZWmGAjS+bytkWckIFHl6/QGb+6TVSXGiqnVU/ykAk+KCpnYo3
SLALHaVaINpmLIHAdhTjGWViGTWIdR0LE0NxPgUWuc9riwFZU7fIWJ+OqlOhYwXme75Tgv6yo9Cs
Ymsscqp/RNdKKftuVw6Maovn0w/BriAtf/lTDJX/sdwb4PrNy8Hhb/nhpAmx47v02SC9mGk7xCq3
vm8ewa++jZ7IbVTC8/5CKBJ89Vem6ETAPTS/79Oj/h8xl8poYIehy2NSE4Pu3vbrum/Gb/AJ43N5
8hyFVjM4j73zK5JVsO3Uyd3spuRW/52H4VKWG1UJZklB/BCx5T/e1aogFTDo/T0TinfuRtvh4nen
hX19tgIDOFirWJxcGsVL/zQVcNEJqQM/wNVo4jz8vd6J1wSRDCOrxazUBV7jOksRW4wFrdJqz9wt
V46HdPGLkpGi9t2Qo+QLwxlgi4bNXb+hSajxOsThwFyJq3/d9HZVGKDax3y8hHsh9v1Ej8e0Lnnt
VuzKCotoB0b0yhd8sPpJYuXcwjVjYqIPSBY6+3sEkerDQicS0JwofmgahvR7UDHBbg2syn5SGz24
M6e5XvsuxHCLDaohVpOPXvmWwTGGTkvI0OhBxEhPXOZe/QPoj8m/cUeE606g/JVEQmBjZfTpLYXo
Oi7MsS/1zjmM2ybadJc6GSF0zc51ENu/73GzZJyQA/3Q3GX8pKLqyGI1LKfxgiKGexKhCQCrE8a2
3oqeGbRa+4AjgGZnRS9O+WiT30XQOJ8xVQchByyZG6JG9JZ83A3kvUTe4HucRGKgnbRrdjtE5XD5
qnPuF4SZE/fwEVSSziLFcPNMiU0briorOp/1SirKhUgNL7tOVD+ehIicZFeLuUkZZk7k3As62Zu+
zKxFROYDhJdGRoVOlWuxfW5uwWzOGhdd+TMdFFoR0DW87JlPv6W/Pc09ps8PGoUdf22fantaRrds
d008NJ8BGvCHtRGvcQIXB41wP1Mh3adoU1ClsdEHxTjkY/bPRN14BGXT78+uOrUa1p6K8qDZzNXZ
ckKuZlVsAJLEcGzoOsPHgz5FG3gUKMLJcsfagTM8+Lz9dNs2121aAXQ21kpovC8vrqRWExmvNxt0
gKxSAYeQfXn8kUVPl0tsll807wwpv05D6znyltp9dprz/ZUYIxAAs3BzKyAJPp7UjkPV2fm/iIw7
zOPD0O/K9i6sl/pcNGzsNlNn9pSIc++EG2lS9OES0ET5lf1RXMPH5Fb1EKKJ4RV2Idt7sT+mLn/u
BvlUAzb7lerfJ5PIE0mnKYFJJB7OwmzeIOhzlqRszC7DIEFOCwbv1ljf7Qr0d1NMO8kI5FJu7xX5
ZROLTCyB+MlZzZCv3FswdaUF4OYkt/e2+ET7lJELFjPf97DYSrrHO+gqyw8z5OZkqOTBwslayk9f
XMaWcOCKegjaeCHgb6PjyMX8j7p42j03S6mkKao7vEVxritKH9Y5KJ041QllSnByCY4W9exvDKvI
02V0xD5iqoRdNd2yramXtHaWsDzKDn5knd6+mhPJx768o4K4euDEwVxV0kBi6sD37TWTF2dEF3ES
rLqTzAmbbYsuFx6+dtxsnVg1wp+f+ftGzNQjjBbIf9q4lTYmnUMACECNePI7NCXZ9SXK1x8Vjxc3
WTCdw9V6i/Vr7hItFX6MmiUcjVFvH70ejCNVsdS8PEuJgEXYdEMQaYBdLf8OG2kU2xx8LCbW9JU4
eqOUQTazQDmRXmx0cwo915NY73kY9TJ6PlnmYuj4sqoUntfkdThk5wyzr60XlFbPxCZOt05hRoAp
1zNxLOGin/OX7fbBfhg89klx648gy5xSC461F3OF8wX85c5WcIdgBJNTuKLMaet4L8fG2EG1WdJG
fWoou3wjk0hMpqyZbOzVP6Jdpj78YwZ0gxiD237reWvW3bxNQW0PSgn7FkHH+LLETj5f1BHM0UoG
SmkQicihwGvpyWFHQX+PMIOnRx8iK3uLqs1z4zqNxFprGNNEI3GGucu6vu+dF+MvhbfOPjD1aGB7
lXZEv1Z5AEpJtcp6XCNYJJHrn7xQWLwkoL1Vx6bU1rD/q0lsaQBRPiejyDA+yLNACayRiv3id1ba
1SSqTw/3L/JhVOgEOny2t6fbu2FQtymJFhVoUYlUgGxafJXCFJUl4nYi6VoJBPui/Ts9EsnQnRtO
2eSABhW1b6iW/6mX0WnEvLzS2Kdy4QqQ1TaG7wuIpr3X+DIQQBSvCYieppY9BAwgV3sRNoZFeB9/
H7gevsTTOUQRCuFmFRdhBozrDz4LVzcTTQw9PxMLaEtIYidn9YzHhJMB1pVmcb5qCuZ4h3sr335T
lSgTrmTvM2mI6DyO4MkSCtWCmDupj3qEzvfpfpaWiwRADwRxyhaFsWxQrR6n9uGwq+4Sp0ILb5D5
MvfVSuloBTnH+iIQzGgEIEMgCrPrfNDnAXAAiHcFLX6a15slb+Zp9LW/cU8L3KnvBhW9/YmncVdj
rvweXxaIQAZLQApIDGXQw8D9dmiZlrrF2ngeapagTKs/v1cuJMyO03cVFGNxs/oYg2K2jNELVmSF
TMgeD0unKAE46K+vDgMMKtAMr/URPQP5xsSj9frlG9NzW1LSYCDolVoic4ifnch5053yzfn1vd9m
LGGhZG13HSgFv3kPAEP7rUSAkcUgX4xB2LjUh3FOD8y16SwdibojI/wovZmUC3pv2adnXcixck5N
uZUwua4NGr6Ecervj+SNo0adXioaUQlxPY15Ry1IGMa7e/Vo5ObOkZO6CxE6mSfuJCMtdTbKtH+h
ieDAvJ4Hxx7pb0i8IEdFXs+YNu5VmVCuewSGLIdtaRnIt2LjZcM7toqiaUdAk2Yvt5MolJVG9eOw
1DzbYGcWbkEh0xOXn0U3cqL+lxzv30xGmhrZI7yCEGITGgQgUfU+sjPlIj+vt3qKo7zhMdbzHugK
+L/tp6sblv4D7NAoS7kVHXcatVNjlrbWkbbp8sG2RtzIn2cdoHUd3LJVGDwr+qEVKhmQH8myGvMF
UU7FktocMjk/uEi1zSp1ofXd9m614Jd9BCITZNjvQ86JuZKyWOS/mNgp8/ZN9wNOjoqHeDdMXAGz
cuc/gjDriGt7sCF+PYpGbnY6FRrDF+c9+2L5yFNh3/Am25aFWCsr0oH8oYBFwBRiuxFoTdo2qLth
dajCUjSDlHF+VGfirBI5j3AB00IjUbG8eX08e4qYj285y1Onm28zFSDVObGJ8oOGdg/UpkAB4s2h
UtBmhYkasLuSRf+5kwWNIWqkjFZdJAu8SzcWW6wiXJDY56KifXnobChNreevm5c/k7+An9SsM1XW
1NSAmV/IfpzYjsXuuleWrZPZSibDzh87LPYXdpNlc88g7iTHgiAgs7NSt3gKV/7Dr4DBov/s1sRz
PPzFSwKZmQ0zjRVZZCrXHoQRHNJcGS+I1OoEylBIOuijh41nCYm/lEfHaly1RRVkAvnRLpRYb1nD
HOQ8z/zcZBLRWoPw1tYRKeyOfHhgRV1QIJmSwxX1EhjR3WidqSqpcz2+0oow2Tpgu9o6HsJFy4lN
Kr46A3vy3VrhG2BOhe3xC6/a4jAz1jX4H7rdTDiqmxmKFHGCJCbKapVeh30RvLLmCfNZ4WBtxWXY
qzcE1O0iOwSmkh9QEYlh+/9B/5q3VN/VvMvi5UzyCWp7E9DFXjvmpr9grcOVRwOWiqVfjX+RfFRG
1Zo60tPm9kIRSY+w4saJievLMdfHyryTPjpjNFFBP8vxhONzCS1njCXF3m8jT7VSIIKAgjNujqpk
A+t32yJuThmLtvVKKtbt+npBBf8EpDqwdQjHhSY+hwqYwBcieDV+uqzQg8hv4KdAONVgLeOV0Hda
6Hvd1E+SBmFSeRqqmMZrWidkrSRSbEU/XsUb6vSA2lKtuqFZKOsJOl3GrR0GLnaAefN1jHlmISRv
YzGtuoMzvSRbMCawssfCvoQltOG3AHUQM4cAn29RtGgGZMxvQSAMBuwvnKAzCX+TRqeOvPfHW6HB
q5lyo1bMqz4iGyeUHN3C3TTuRv5ABeEWi8lABL0VDnj9tchBJP0Z/Va4Y9AY7ou9fD/NHI+N6zxm
GmG+w4IzwnaYzqg+aHOujl3mp2eqJVQOiL1rKBh5rPWIsXfQb+YWXKmH7k0WpdlUm62HvVQTlw9Q
/pnwBxCJKJIYOITfkdDmuJu4sNQz94VXqDvJpwMIOlaosK9S4Ninww5PH0tUEhNv93r3HDJZMXyR
6E1nFG5qKpyF7VPvXWCtX7SGtbHcxsa//akQlXsHum/hWrHZuiOuWR+fhko0Wghtau6iPyyrPKPD
k0M7jFOsctTl7uGuG86CfqlaoePwI6FM240q5zHKaSRojbDotHHFhw/1hTskBvlIs3WGZBvwl0+9
CPxUeGi0WRtOxI8rpFx0E/KFcaDCJWz5pYIjbubCcK0eHbpUn/AXDBUfOIjD+HNk9ECiNWeM5yzS
7OETk8sl2C6nenQ4KtoVlG+l0yzPF1xfPegz++QE3wyYC2ueqdaJLlMUDbD7u3sj7WDz9U7DNZiL
ljB7r1Ib7DvWpLDuBEPSJJwsvKMVI2thxSPqUlCxTl4kmJsgjEToF7Xi9Srh6v7BobXTdrsim5Of
GSWdCzcG59fViTn0/kiUhODG7hNPfabL4fSiq8KSN2Eynzj9HT8mODk0J6OHxodh0ESHG+kdT3zr
ihn4q3o7MxSM7JLS67sPV6h/kJgA4GLH77IgNiswy1kAwIkfIs52JYRjAJzZ/2yxLIehzaXHqdyu
FmmtO3MD9jwzhgf2OuZrBrSufVsjwhIM0Tn+zhlDSA2gz9yhb+7t46npWYFdFgh/PIyTIAQaR8cj
edN7oenMeq32+sc7tXtLyalH7GKGSYoy5nJqLd1bT1Jc1KfvVG3QJjkw08jxkIzNQ0lrdB+r17pQ
FZdfrrke+8fC/M2I6khgpe+udY8FZPeDX+I96HHFCvNFXTlg3EWgpZUPX1juvlU15ugflstvqEWM
nFZ/ctWUWYhVXLxpeBAK3G6Q6i0wM776N1gBlA2qgoUjzxhC0tes7AfShrfnICjcvSnQW3Zq1ZlM
wkNU3vKT4FX1tjj9ZDzSWZH77+46sca1iiZVj2kamyQOzKhjMnDAXq2HDFvtxuLVqPmrxH3EH3qo
8PUvCgaTi+Oq3gD/lNWXlZqhbuvvPXNVt62bimSuO2ZpBflmAbQ7nW2MLpiJtzsIP+XLeN1X2sV3
NkhDnPqy+M7uGFtr65DdpBNevkjRYQEdw+N//iHGRzSyGxTVheGfuMQCjMNmi+THRV9QrK9gSj6C
5KHNglXOww4Z6jjBpb544kZal62ZMbMxkfqMx9dEeMW+WwTE0E75MFE87EJDJD4mFn11QZp6wJej
KVEuK36GQiTaFgjKMHJeze9zibteZ00VB+QRnrnb4wEYWZX5VPOhjl8Tkjamfvykgv+n2eC/ZnKK
EwmAAdT0WIXctv0jgKPs9AYzPo3WZ59bMtdVxUj9WXfWkOIYiHP+D73FhDaoJ7YPedL3wXsQBaP5
YQbDH5D8orN5171+9cCJ4HGTFfHiM9I3Eony1moWsrc07OtyqWKIUuhaR7uoVm5cRP/oxpO2V5KF
Q3RwSTDIVl9Q6IRfKkJPHQ8npRN7nEq3mUchwUNgDnCt14ZbFkPDUwl5ACSR9nsbaTnZHGD9C0+T
xGZnYfFoquNEkPo5tfBR893HMeLkRqP9PqpX+f+69yA2ziTPhbdE/G2KF3VYIPlUtoUVxoY9XDQr
3g7OIxc/m3fkEuGV0c2vVn0TuQkknG0JWW9UzTcqa49hYDYB8Tfmgn2AEZJbRS0YmRR7FrzXkulF
hQnY8kAGThR/DjEWrsIRayw0Yi+i+36KTM1fWlpvB7EpJaNmHMKRf+yvTgK6WO04VaF/W9vT91un
7iPud7sAGYJUWEa+qf4Dwcw9G+///NR+EieLbvInRtMePo0dErSVC/ihVHJare/LhndR7p18x2mx
JqM+/BaV4nLqN9trh8/YXx3md4sQKOhSzVw8gopTgmJwGN+nx/YC3ZSn3k0jr21onDQ08M0vAixz
I5M9hdVLPPoVwOoxtN1+q/akkgvfmhl4lOViwudmu0+PFP1mwGgmQxCF+16WOy71ihVedtuZVp9J
efPeewz3hWWigqy5d1+q+awjdv6HMs2owN3S5dJHhVcC2VG35ijX5JejQ4bVN366hbicgT/uR+oB
TORbbRbb6+TBMPNoV2cHdb6BMZr6rY7xRwH7qbapWvmIRs62hCgpLZw/YWLE8UUsLAe1eJSlgraU
mCkF12cjIuuXJFV1ouPVEwmk/lSx76IwfP4Xd9hXDQaYs6nh2ywhSJImUTKM/1l3HL2JL4I4QWEr
lkXmV3MgVpsMKHoSDKq1p5dArdUW6OBlY7gT8t/SI9Up64tmRM4c8kmlveR6PBjdrl+1/UlfE1CF
2+w/yaMcgtNddMQdlcxfCxCnI1nvuOODBWpqV6ujsjJvs8Qw6fTUQBVWZTs1ju5UDHHAVWCXG1Eu
AY48ZbYAS7ZSTzPrJh02szWV8xq1HhilozDBEiRULngYIxvrhVIEeQoKUYe6G1T1+w6+YYFJm1VY
7RdXy/MfKXLLN7U3b2jPJYL9cxbn4obbfaoc4aFQ5wQdUUBfS/ALUBlEzGSdS9qMk8IEDnTAv8gi
jV44n+dWIP6J29PCoJb7kFzPmq2AAFNddr7LlZ806NTr3756KiHU0hSVF28Z6Xa58GnBZoQ/Wbvc
do/vDSKkbw36ywQQN5BPV6kcKBTUMLDiqxA0mJqHTc0+5S0xGsYp5i7XRtz32qzzxGGu+xqLhspF
zm4z8YBsaOlyr7n+cI60Op7UyqhsqwkfjSgR19XdZx9H3QrLEqUrWjujO6GEe0OJUtoqFBD2JIbf
kzTuJLxtKWkhZtluEOM+r16ffnt8bSdg2MB2ZWGzBLiaiB13W1phfVpI93uBzNnR8lPA6dfOEp2o
brP5wXRm9qKhqYnt+p7WyJYnue3If5xCo4qgjCiVHHe/Np6ylV+CTofknb1UTDnXs/nFZmpcJ4aW
dLEL0+khfE5dh+70YAu9b5XKNdmxksLVrk1QsPNhGSdNG2IXWnVeYQI1YfFU8FtLswyAiTE2+Fk0
rEAkEeQJeUTFBCDv0SyYgxzUtsSBiEPLni8nPX7/FxpVW6yJklPW80v3ytH+KzDLcN0sEQwEz+O2
7AhDCtPKqiOxUtCNZejSU5hfCYRouRUb6GpmzlWHrhQIyIIFwVpSjq64mKzlRrHKuVdYoqTtNYIn
x+aMGHHnD+kTF1Btd4+U7amoDvIiURc04c7YZx07Rjp1j6/JYG0UkXp5MfDyv0nNUO53iqDEDBQK
VJM3NwUNc7g92x1vgTnutx40ijfOyzDGNH29NaEg9HyNkwKUKoZzvgno//PcQjonbLBfXYxxwdPY
kAOnBItVAQQljEpM8aaEcZveAGPBSYldHcV7/BPxfKBf2TZ4+AxRClJjIyQyfTehMp9GUjwz7GiM
3yKH8+ZG6uUcitF+8mBMqqVPumQa5pVfSpul+C70pQQFHTXJrrL0IzHINl29WgaBgJSdUmpeXybw
dlKHyMsEV/rWnB8fAmLa4zaz2HrFBp0ZgejproMITXgz78JqlA4CI/MDaV56BaQatP5SRddFM+j+
iGdWXQPBTyENr/9mbsDb9u93F7NyJf/Ge2181GD+eMZro2B9/NTQxB4AOY859AuZLBXYi4/Rc6+1
R4wvF1/zGOkYWNtwQ+mSld1gls69M7Gb4iU2875EuB6HllUjYh+ZkHM3ln5SdgT1uflh5UZR30z4
k6I8egyb/n0sqjyG3PIoz34NoZrs6FWigWO3ol0zBF7aThPe94WI5hUb0aXzq22d97R0R85snu6I
mNisT3o3lz/Otg1Pe/9iIdMiIbVTm8IGdU/ZkIcWjkJqI2BIb7llX4y9XJ7aWE/MORFee5YLEEI+
UcsXm+O/lYbkJ18zFV5gzmToj4PkCuIJ58+ce7Yviuws7cXgkX9SRKg33tpGm0W8uLqMsnNjkzka
mguXFSbPSI3auMnsRmcaWafZ2l5CFfu3BNp/qTUK49Sfy3Jijjo6qEBWUszcFSdWlQDuPV1Hc/F+
encijzDQM7fTMUMmJK1zB0fdiDGcG/6Bx6Nz1mN9YRveyKxo+Mki6BE7c63YjMuGL5gawwT/bs3k
TdUt0yMhbEnnxl9kodE9bT5AVEleAyB7y7aDwEQ0pH8P38Aobwg2w9bH8F0Bcef7fDnj/zesFt13
ivvVexglmBzpyq5r/mRV1qjAYFmdeegFYFrzzQ16/YUSXpifyYyv68ikWAuKle6+YGCV6f2r5dpb
l0mpd9XDsg6Uoco1hcHDBjNvgHLXMl0Cy+nuA0Bpxe6oo7FCuLR601quSRfH13ANrcwtBUDtT+b3
4x+l2u9p4vcWvd8301svDQ+WRGcrMGLKOk4ukTOob2Z2qcMHFoKtWhRVF7c7PQIjmlEY2HT9jqds
OPfXuFvCwFsQC3gS3wGzp+fOBAjxTYPR/glCE+azjsTCWtk8FoqDUfYLg+Fp5GUDP3Rtv3RP7NeF
lACW+ky2504BODYtPp5YJQFESlw3r0JBjCKpirTWg3JRgo5YHu9GQPTBb2gz1X5Ai8xuiz6fPSFG
IoVeMpdOQUseNPaHatg6bdHcvAFwG5sQ0lC0mQzXOmYoS//P1V7tuvS0K8e48hlv/cqHCZN44ojF
Xic0kS+iKTmG4SzaoenGNV6/DVENOYWENlEYCF3Duh7ssSeK4jiRlIl1atsu3bq7VlqN8xkRiSQX
GQfgwZNOMgRlpy4o3Cibat8s9ZC6dXBRlOaFL5NKu2fVEo74AX9LaIQ8Dinl5id4lVdjdywZgEQu
0IVi8fdbIEvbCwTq4Uk/l5TH2pAAjNSSW94f33fKuOlqRVNu/ZXWoAr122kpJgaziBRYd4+AdKdp
FgSi3pfPr8K/zLvGMlfJ7VHlNxDl4w2TC1hUw7ieJtudi2w8zex5+aGf1kv6zBJyI/cVJ2kMVxBa
OqGXdZ+8Vx6VCSc0LMa3qRSE2AKFNQNpsuEz0h+XtI+1GZQIiW7mGv4IPw8/SgwexGZSwOUJd9VH
+e2aIDdr3OZNGFD+NkDsh0ENS04qWRipzp0Z3AWmQwdr1U9TJu8UDcVX4mezj/zNdPuS0AQD4SSI
Ezv4IGhHvTk4OOJGp9Wplq1lo/wj/4C0iCSGm6s5HOioxDl4oLQZha2WCWvMn3fgzx+vDMQ0DuC6
ssO/bG8GRjQcFNDlE3vea+O4DEV8rmSHPPZY/JpBh9Iqm9gQSCYWHdaNmoC3kn+Fg//v2ZoLcQcM
SsPfhvoNG6FbCco0mgFCcbTU38b8nDGAjGFYaypbDu0EuJXYaIqtP27Om4N7FFMdAWL/jH7GK7vq
cYNlzstAjrbIYAx8sv5LfpQK+3ie7Je663U52t95L79X68lp6cM+Ai4PHbZaA6PaE/cOnv7AjKbf
jQ1en28LpmduRLG0yTiG92Soh3Pw2N5DCGMjVLN8X+jWZTjnjacpZeAkj8UZcdvvIsMcZLJLhE2B
+KsfyumzD9YqgXuB69leLoSfzmGTADkKhKYOk4oxL/NgTUuOX8wWQhs8fsQIJFbgbZbpJ9sxpHDi
LQZFkSu2N+raJLoFiRZ7/WoWAv4ckZjO8Nzgui9NemDEV5aaeT2K6Vd2KZtfO49yUmcS2yn7NEhD
4+eROrI/Mm6T9fHBrvMB8S1haNVi4sBzdoF8K72D8uN35+foQkI5MdsRBvb1dgDEXhYwKiiRux5W
gTn09j/0lbKTJz4UZ5JwsDvR/vkhoKo9BJKjIL9W0R1XUOOcV4hliEvLIVVT+Qgm6PCzJq72irU/
7vnRvakYN/kNozyGKKf7TGi6Vd/fcw3BNMjs37rCiE2BvxGLiBsyB0XgS+/sN96slF3fDDVzvGaV
41r1nMMJzlB7o1WTvnFmJOgTXYBgLSGhOVU1aq2fWFuez1dCkVJI3oqsXGJB/R6iPTwTgqGvJGdw
K4yiuTttEpEa4N7qLAcI4uQI41SKkSwH+C2AiE9zA5D4wzzoERt0hhf5MxmMwyXBnsjaGSoB36hj
zIfKOef8cHjDxAaX3kXlrnzumnD0WYguQBv2tjML7JmQkImIq02fYhDMCTBhoNnh/oIULjLVBrUR
tS67tUxsrGylzUnhotkoE97MPkOrSDv6AEclCBodjbnGhbRdkk9VTjTvJlWe93AEwNauD4rimqEa
VwCtlQryxFI1bhIokn8SSn9vudDRe+R3CuNsTT0T1jgZOUGSxsW1v+8rSYwrcuv7HyqdL2N7/MWK
kpqxp0fNFUQD4VNVtCPVQFyR9lnjUdSnQMWz7UsWShlCETmmpimN6E0xWgi1QP206L4isl/YCbqc
75/U3Gct8WNVsgiP4SCy6nbiqRCs4bpNPHYordAYAZj3YifHyTIO66/8KI44cNVx/yeSqeRhsvZx
EGIcRY15POa7q++3WwVur21KxUPqUMpIjQFS7YW/uNuNQt82erUN0SalkfV1vskoAwR7vRKdJbT7
+GqNvaBUw56goHgTTaqEQAPT9KeXivf9g9BYeKSSae06BFh4FPM1rc4Hjf47AghX/XsAAXoqifnK
4ygShDYoof2m6ryTMb6FzoWHmJKwZ1VSLy7xvZccpcbjQolwi1e93vdtkor1oJtdHN7Kjwcln+0+
STBSSPDYc+CNjxDRnEodigERgdrtTSaY0FgEWVLyKs4YGsfopwDgCpddSxg4Fc9eBjb3oTILUP89
vlgcLVHZwtFJedhnuf9eQVXzpzE4KNh5p+NcGVoP5WYxIhGic/XejfM/Pr64KVJMu0TaJBISVq7E
cEF++EJlLoQg0d0f0Oyn/hZQhQmu+UzbMbO4Fm4/EJ5pj186I8BjK8MgUQvd8Xb8hI925kAwJ7ke
A10Tn8i10Q0eJ5SIbY+KdCAs0LfMnWUU5pQfOCUlK2r5ywpMX0DrEwm9+8CShtndnYk26yVzhjh/
vHZVlbJiHg4zt8iF8Oar33Lj3Gjt1+AWSd9mYlqMzqsUnyh+VSuYD9RvW3/ZO1S8mCUDuST4S3BJ
3rlPyEKxmAEAa/qxbr9gXmfaqfYJhHAAoD/6Qi/51WvS6WI7ZNR6J4hnM2J/JPAXsAiuhBVnsBYT
AB8eDl6s6AvutqEWU5f2B1+JiAGH/9ahZFXA6z8AzemjEZNYkBsah5ULRi8c4+wxwaYeSJYaK4U5
08qAmwX2MkCa4d41cktvO43d8J+3Lwcol1pLKe7xFakhpIjpzi32or1+OawGhFHM++18V/UtF2Li
NM2+FIxlnNvePPZUfTAwwqjQiDKedAHwvbUzlpgTOIyEIH2scS5M65QXnGb5RBUzSdgnUUJiDy5l
gR3xVoETzS+auJCb5mV3GhHuoTDFeIzhQnvWbAtMy2niIjvNX3cidr2Fr5Uh5COSW8AHdJq0zjGC
qa+pc4UWm7i2MKnOiJugo5dl5D8/x7LRszr9PV6yVqXSH1YRnKOSS35w5sz8sqxtRU1Ke1he2nLA
ajPW8+PMb6b96SAqpvy0xwQSFLrvW9UQXSWaUxyWbAe+a+Jv5DEmsv33eqwuUXfxgmvu01ZcB6X5
yj1p1fesEiJMegQ1gK3ALZ0VDdBhPcfVrJ0FGNQQ5I1/Rk0QrvnfxS092ftax0MMU9yLP/HvtEL0
IrOOfG0//WrDm/AJDb0MpLH3jN0ffU0xn0xQT1dGNarDd8llTu9r/nbF1jBuhW7Cm7zCNNeHjTjm
4Ygf4Qu5tu7Dx/A6DLN03UQXaRBxBFZ/rIBa7DggUE2HLMaMm7iNMayuyaMNDn1BAOqEto+ahk+j
kl/QCX4gWoG/Mm9c1kptjNllpurBIZgE7bQ8ysYfDYpU7FMjLBCkSLtqcCgiZE+xitcaolZmfWFU
BqnWUJBQduq1pXJlAWoF+PwqZ+ixarMArodKGUD5Gog/Z108B30V+Y7Ni5BmGkuY6T9JMQjnsPXu
x8GbjK/tZVuZCfi5nzFXfXWP/j0M+A+zsoZ8d5+ebnSc5k3cpoNvsaxZ3V8cdfzh2aLpQLM32JnE
wZmiG2WYzJAG5b+oI2TYnrz7GV7715gV3QTLFrPK2j3mZeYYLyjT5dlLDzTjarAzHNQnFGJZ+Jat
JOBWc+7HsxO0X7cb4MK2NdeQCtswbRPHqD6zG+ly/Lz3WS7Jl8O0D+I2nWPmd0HmCI52CBsZdt8R
2lZwq9L7TSliGCs9P/I+bzjec/a0l10oxw63BumGJwfYX2Z4ftdSTSl9fWox018774EukOFKdZMS
mNzAM7vReAqjVW4uDZHx6GqMan6PqZrMg5G3+A0N2djKPEl823WojkL6rM6SQBr5KA2GYbquJ48Q
9DA7YlHovInXHfvgRqSR6KvvVnZivE22Dh6f5vfte42B2TWyCLttp7C2TRTTS7Qnd+I7eQLNaulr
h8zH7gBik8BlwfPhPVzLLolcc+KIVEfhNhgL9C0hc6NEfGMU4mZqz/kfSx7lVIh3ushZOywfSzr3
atGGQfub5b6K/pXBHZ5LTN7BWiExHPYyT0i+ep9YgOmQWTOFpUa4ojTiNkzG3LGwk6tQrSncBIAJ
qEp28n1lMQn08Qj2RCUBJixxSttXsby1IIfesYAy1/3S0pOsHBGrpw3G3N4vp/xdd5eQimwNWCpQ
2vgUxZnx7yDuxyrDQmjPH0XgQxwwF/eLJkSvPqe4zX2UmCnx9tM+rg9abgp4+Yhw8CJujC6kOlVX
GmVqqqAkngI+F8yJH73LoBW6zjrsPd5vjzgAbA5FPemmEIZ8k7zRIexZ1sSyt6f4yMcMAj30UN6O
5CiqNTD4PVu6zTds9hW8qsFFj2VCu0cgVkPinF3X+1d/pCgGwGKW+/wk9lOaaG0jK7hNhFtDxNfI
IPLPjM3mtZ8cR18ZbUCjid82yYyY/Dd0cGxR6Sa/98Pq2OyNB+fdcBOx2vUYutSvTa3JCQg4XuEf
l/kxDJm8LCoY6Fkt4tAQ9l5LlUFX2UVc4lTUzDS+0swAfXR3avUpY9sOel53YYQmYoikTDdgK00l
RBpL0sWsqQ9yq2NKWk6/mpYls67zM3ZMeQUUcteq53kWduxGqa5wRJUSNf32lHyr18kgAst+Ih+6
ouDccsjXgv0eytiMwv5LKnAfFjlASIJU8WoCoy5UgHEO5ZobcDpmtC8trbd9BCILxcYX0Zkq+9AJ
844dl7OQjbtFhOiw0OMfbsZX28zfOQDLNN3eywwp3qJUa3kEkqR/P+c2MHLuw7pxb7yzLZuP2X1R
OtG4uFOpW4xkHdZifh78JXAkpUymBnsdfFzeL3sHsEcM5gm2ouHFJJJrPhYVs9pGjfaxpjrQcUzN
KMFaHuhStjaQi5UMRw4nsQMEcD9cxDELB4GFSQu3BPXz2PHEFjRGbQEpGAZ/HlPliNhgP3Wvv0CX
5pbYcct1W5TrzvYBHmXSQJo35i5a5rwBIGniXOIFulr9eVAhfJMum4nv6mj0arOUFLaa0jjesS4j
hf2qwo3t/r6smInveI5yMw2Ao8sJ3slA7MmKVUSHpxPHoUZwyUt+RpQtgOFJdqv9oAvSwBMhWpCR
XvVB1Rp/x5TgqDWg/yGCrxh0pvs34Gu/EMw2o+5FFVzfrfkhoJ3QJ1F5LDC8qmg+ytGv6RqhrIAM
NEjrm4YFP8TPmvewvj/kfPONXfs9wc6EMdK+/RVpdNBUow5pqShLvz9IlDx2TapE+qryi4M/L1dC
k6oWDFXhOtBdn+iMOhMWI8v8CYDN/ttaPZlSeINZ1M7BWKankXwI07P8jPqbHsm8Yrn+SmChvat9
ubdYRW786EdhoB7t96oV7pZYUpUq2m1ZRaUwsljr1A1487VZJkhLUxNhQI3ozSiQTr92ObaKCLaf
yAFngzHVz8rucNXkVOt8Rcn6TH01bm5MFeT6kl9zdiBFe0t3lSkYXRpl0D/GLAiOdBo24sdcTGeX
6vFQTKl5+/kHpZEr0D9qgCukerEQUEbGjfznrC6vtWBXfHX2+qqMCPzdHXc/RHRwaQwoQsEO1MZl
G3uL64O2AOOhrE3Uc3L5ANDHPK+0H0SBTTnWy++YMFsSRT8GKLJS8ZOcLfY+YZqosV01EBgBX3OL
7Q4AcKD3NoyR6JczYpn3fvxyZ7FAb5hKouVLGr5gHHDB+jvuoE58/RJAn8OgQ+UMP/Pld2k8WBeB
R84iWQ/BEDc8E9CjhBRJUjZWmfsnsCwlaXqJEJ+2mu2zDe3LhlFSy6ksBC5Gfs1/s++YGyAT7NbV
KzYncXIM4NJIHB08M24RhCrLAD+pj7/aKDnsap/Thx9qW9Q+qZtWdvurzfnLZz9FYlJKZNHDVtdK
USsVvceQsU4Pd2SvMZP+H5Zc9FQ57D4gj+T4gNctZbh4n+jFNT0cMORo73EKfy9mFrw9L2XV2ZGZ
7BY09vAEVXzOsiyfhwPWDtwp+WjCNVFznbCTOnk/secxaGgX6HUL8aMF9SkO9BSKFQpbvIveljZe
EuFEPeSmyEDRW7uRlZ3eh36SHvafa+KjCUt6kn9X+5BN//8JTnJhBRV2XcwJ+97F5WzmWx+hNwAS
dNZckf+pZiZ0uu8INKYu7t6MHo8Ez1DbMaOHvn6uLjO4NBwkyd0kqbQAe2uXbntB9i8q/j/fMS0W
9M4JpDTyV8vj+83RGklvudfGQoaT75i2Ji/oUDolfnisb646RWGshPj8hFu5lvlbKqtkbCIo2CQV
A5Xe+4EBja6ksHzjskmuVSsWsUP3W/LLnXBHWzYP0VD38V5tPjZb6I54HsxivCRMA1isrl/9+GNk
fx8QJHyZEJ16Q6/gVMov4kI+jmVcsukQZcnKpMSrbo4hiRoDxZqXMxvQbYj2BEwmwplLJ6nBHscH
7NdWJ+yr6PX5zLD/oKfV2VZws5Lbm4XxeMOWBVwEJ1zBUKx5JZtBkABik1ozMXNzkvUIyXLjauAL
Uxnc1d5XwrhJMDF5fRkrStBLCc+ZjKUNOqmpCYFrQu+73aou6IjZP1aRWANLoYo7hpK31F6+dWMo
Az2FNqb1XBYa2e0ueNyB56/ZB/cELUQqb0zhW7fE/uFPejWMpwYJZC6l3EkZWxy3i6eLnWe4fLhL
9/b5UrOBklwTmad0yWYaNYXQtazGKreotbB3qbhmv/IAq7UG9ziwxrMygvhtjEv9pQLyyvg9oCei
LG8mhEbXxEi53k3Ma/iKQBGIwOlFkNSSRKU7DAVDLVixfJ4/4YUr8T93GK/f3liVgxH49BAot2AY
8L4kC098/FWBCvVTyGGw9pa5URhyfnYs5hA81lPlyPd+RmzCv8wt5ADha1o8ENZLTvyfGlfnFjGZ
bQFmKeVqc8z+2LSkutAFMJi9+ULBvvGbhCaV6zQhapoMzztDsiCqeaOFSIn14EpTNe/zMv9FQ2LQ
N7xqIXf02CHg/iy4qq0FgkJZawexCgZlW60QobKYwV1z77d0muR5db9LvJDd9KzukYLtdh6jdktk
rYVyEgvKc3CaPIxhmKhpKFK+g5iBMnoIXlv41J8JF7pMmJbt0S/dy8hs5AH5ZJa7Yeq3a2dVxnEx
x0PT4q/I2e7mFgGzwgj8hO3D0C9O0L89QjVY4iQ8MIjiKsMnR+D+gxCZtUf0lOSs8z8anz9qGpjD
KgP8DefDC2YMZ7ug6nCyBTH+bLJsTdBx8rjO1ltfOx9U6x6suH83cV8agfnPf1lYzAMV3lC8Jnva
5G1EDNEthJZA1Nh2O4/neVpzYFbfiJm1VwMH6yYV/+PpzXs3/XSSFWTNEy4Y3SSQ+czTZupC76gA
09ERopFELsEbzlxHkHvIh8Lbf/p6gUPoRfhgoDv9XKUfAoJ8Lcyi9QyVw9h+k6sNQgXDX7PqFWZl
QIJqe8WcpFvXLdZ1zi91KLhkMf0QwRsl2MhzXiX8/CAD8BRpYcmmxaHE+BfDk2HqS87xuWR6SAbS
F1HSn4KKQUnQxa7yfbxSsTHVF1xcX5Ry51uLCfGKXM0YZs+aFk5YZ0Izju8TbTSmudVtoBjJy85B
Q5MzRixJqZQpeU35hotTaE43NbTCrjkbyWOsxX3co2PlPJVeUBg/3MkB21s0bNWMszPAFPxE92eA
c547IoWmMTwD7hZwDD6Sp+NQuKOfLv3vyKfSy0CW9Dh1Y9i1JR1y/3I5bObAQ/EyWLdtT0dhQVgV
y7uaVqePP6FKQkMyesQiIce61k/Vx+6yUZhFW709ZkUIdN5Sjtuzkgdij1rZQ8kmWQD1nHD7kchu
Hrsx6ajZXuUXCiD5aSz3fWwKAG63Hk+e71DDjySmXRRg0nFrnNIOmtXDYAqGKkfM2PBEM7/ref8m
Jb8PhKnIZf8nxRSTm8dQPDv40vw98rD+DTjvXTkQ4pSkFv/RgLT6ydNjmE2L+aogHZmq1zXiCqJa
DPKCe+WpnC2TcGs2kKuS0UYYD8LXEcpcEqor56mHIfxyAJxIS24W72cVjkjTJ0Hm3dY4gfK61v9m
IRPbez0BSE6MSeCfyqePa0ibKxCJaY/b6iipPxNPdnCiUV4VNW497tSqNqtg++OjORwifiX8jebz
OCY7YvelW82pWSpz9B6J+IhDkwtyHzyHP7yQV+NOVgMOhHudTVs6SzCSSWiM3NBv5TVW/tZcIoaC
ZprdJISZ93/ujAjSBdEglpU6EMh8ZpFOcDGu2Sw5peqWQVS5wWdvxCxXRQnFZaNtxgFRw8EnQ12b
17SBGJPK5kppMYlLPz0pf4kdaQRDCeXQ3ZgJEulkZqgNulvxYMIwvv8Ez9Y441BxLPGkb5+jOqbc
tehI54hA2EUK5o5tiz3pXc33IpvCQWcyDfTSvz5wt3tqqpWjpOr0BF4NAA5n5nCeqKKOhFUYUCyy
7ktlINOW0t5epaK84SKExi2i+tWOSTynKFFxQJOLDhcvOPa6Mim/oGhKalI1VxcsS2z7Ib5TjEuF
uhlnvtX5Y1+5mGnZB0t9I+fixL8I+fI4AqTeT7f+5rn/aNE5Lrwldf/F31UB6mAf9KozV96WaGAT
Nsw9LRsxcO9itcE2W0i0i6+JRFPvLZovrSEPklIxruwULrYMGqHsnBSx45bdCvglqQ5QZjm925z5
YxyyBdgqTnbNI3ON+qZYUI7+OeUfYToe4Kfa+c9Ip9ntjaiaIhhtDXUrw10uhRg7uwn2FJfDXiL+
qUPTdZEO76X2sE55idQpV2OpfBushLC14PeUgnmLjjKw6mgM/dkX65U1majyASpgABybeanUyZ4/
TroSzXkwxqNB+E2blVspKWrBA/eIlBfYxl/gSNmzLDoV+L5cddT7mzaQhEyZKM5dQSnSQ00H7CdR
E/wmM/t65sloilC/2EUxhYlfOToLChVZQY0UQOCVRb4uAzhKvnAweStkvCgZjzLT7UFtLIR/R2MW
AnCNLiXdEKEtX57Ykdvzy3p2EEMt64Hv7kL52dv/ptSTEUbrm9v5YBeA+Xr4PrE7SXq7MVMcztWR
sG3i7BN1b143o31sHdYW9H6CSVp/A/JbFQGW81Ma+SNq92xA9wVTyfx15BKNVzVgPPuqmXNJvO2S
BFa8PTvMcbfaf1mwgS/3npExB3X8jNCWluB764ySUifQHTmx3/3DV6LSBA6ACyaDyj6YpOXpVYjR
5k4Yww0J/GaQD0p9q5iEtlukp18afIUh59teqgTbsgGcnEgRd/so9iIdWPwPLKaDIXD5H+GZ/UYu
cf+aCCAO7XCozkN8I2pxP5vpdq9D/QOgmcnsMGRFj6h2b08tCeSv/5/uvcvTy5kXKPtsjkgIRysK
A2/6H9QgOtFw1uqsmyO3ThGTC4sgNZA14WxSTW32XRrZBoy/S6zA0ImRhG2lUQ9Nr0PB2NeqsCaY
kDc8yb/l1bOd8ovBFXYpXCmE6AkrR2zn6oFfBj5PWXrk7oYNg1kBhM0f7Yy9vgrhfZP4ZbDNjBi0
jdEWByl6w19/pnA7lRofelJwjPL1QRk7MAGPILR3nQj79gUGpKZv5eUdxqcw0T0yLhD3tOwB8eg1
mMSQuy6xGFeU3OfRI2nU8bwtZPRmRaUypCnkZWzS6gYr9v9/9E8RJbGUkYPXHy8J1OkhKJ7KPs1G
CaBYS+SfD2tUt9PA8vf61XIZbW9+p1MeHHT+yJWmjON4x8vMuU+9KaMQIw+JaHDplf+nDl+8W46o
YzyX7zsV/d7d+SKVXUpj4c/HRqXE9zo572iqXG2e2jY1Q4Guq2owiEwrEri/aLjB9YZOrwJSZ+fx
FzG1JowFzo+wZtO0EeeH5EfHn6l+ctpwadE2q92wFiAifde09zSIsaVBjA1sdv7hS8q/dpp9ruiB
1QMy8F9v09KqW8Xz2rQ9hw+9eOSbuPkX5zmB42uKka4LXZMrQvKBkCeGp6uZWjvSaPBLT6Xyqfhy
scYyC9S6FjozpC8joW4W41pSmsPM4DuejBjwz9/i2Pchb3fijdlmGbFfUy5syET7qhDNk7E6iAe8
AjY84V/1lfoy6wROAdBkWSbLcnEw/w+V15G4EKYV4JRGNzhiqq56uZShUcr2Ga00naaXMHn2Sflk
JK2IoXFw1TdOP4Z+GXMrwhYnkNIBNZ4Iva4oJ1c8xBAyu6w/x1Kh8g7nvWM0FGK/N6SWim8e34tH
uKrTVZ3gNOO1VvHL8XfZ4SJ7heo++W17o8W4N/BaYXN0vaFnh9XTR9ze4U34dWhUAIO1coR2iIF8
qFo21fDuubKB7U5XQqD/H4QJtju8GBsxj0UeDYNElGbmbf3bRNGEvMOtvDjO7gprpp4gUWgda482
GRl3p/ZXUuuti7mTizIdnN9mREbzj/VVxDbmCIQtKmkpbzvpyCFZ/+Mlj24Srhkj4TRLOslAB1K3
h5bDGWp4moYMUOPgaPZL6+0tahTJOTNnrg6VJR8ic56eRPT52Jl77C2QGZvbtrGhTPN0n4c18O3d
Nu06gF3ZWXwV0/GGrUyZu7NAga0/CtbgR5yy5OxID/dqiEQVRRqh1So5cWfmglJ+Z6WKoOti3ptr
sWLwrUgdcVke+6UyzRdFWda90wsiNZsukHKPnIP0nDph289XpD9NFYlC+/cRX+XI0MfpbuYiewV5
qH3hJSeZzrYQBVB/S/FeKdSoe7C658hbn8T0MNa0WUChJkDU8hr+xIe+FdFAwULLHyA/CHsvF6JJ
4ZQTQw7nh8J1rlxA4LD44aLrqdJJYgtAIXjRiyuk81nMvUFFRRDIzHFq6Epu1RNwh06+QSzpqtoC
ORfAbqFxoZYydTAh5PoIus7q5l3Ra6/XE6Akx+0SiXrIE7+xi2UGJKqehTAxa/WTWD3n1LfzkC1N
5sHkzfODOQqI03w2JJX0W++M51ib3lugdjVHuEnI4Wx1g4+5lj+TjyjAd5R2CZH72KbMk/OpVhFZ
9O5+nk/gQLw4tjSOfBR/gK79oNABIABUAVzWAX6HCyaIenFb9mD9y/emdjqvylf5RVnWiKxKp2WD
lhXn9gNbwxl61W6xJhTR7EpCBS4sdue7BiiP/Pe2iUz2UJeG6chdLu1In9BlsOQk4haTvXEmgCF1
gFMsD5wjcWGtClYjZ2TP6n61MzfnMluik1WRPdoaDzLyK+4oRwYVaGhIVkB5ovcWBdJr4m7C8/JM
gwOlNgbY2fq+hq47yYaWM/Q3GP6IVTxCzok9hzW/np/JNgepZWG30vQOMdA8HhV0NuGik0ylvrzN
bzofFE6Cj/ZKR8qsO+UgLLLvbt4xiJvF5SCDf5ft6PByjtWJbikn8lqC6a7NLxpqO71nBgW9Wog3
Wjg66BidsmcJeQiBVMPk3/SUiIJJTmrPbuFJunfGa4lRALN6TgUAM0nQGOHqTwXY6vMh57o1B3mK
6AdeUJuBjqLW2Zi0AvHW2AuIq56RU4J7e/PXGHvABnAV/Kvdgs9/9crv7+pvQwPZLnYrWwDo5Bc1
CMMhKlJR0ftJTxCOgwqdLZoLJZlJvsaoTIzrJ6mXY2YHqDccrXlmb3CQ0qzT8PjemgRzxmDsUArt
uN1gIxxB6qFSBKkBr2kx1buiAyXTjNjGQ4r+2dRnIKPqnBtX27m2CMG5jVDcHQmsZmcz58mhV+Gy
l21V1EtnPzKH59k2rVwT7RtHJhpE5qJJbGWnftLhzPvDh8tEBW5dbtJiY5HJY/jgx0DXIFsgsizH
GmrF/TwArfEOnUMoGSLDJNgu4099fnuqpYRjYfZVdqCt35jQjIDzF4/OW5DvPjdxyCkQkzjnrNY/
A1eKszU3haA7NbPvXRXF8q3hVLlIys9rQavhoDN2kqfaTkL8ncYZ7PEvXB15XaHReJrxWu3bnB9y
FEck2jS4TsVa/f+cFh+VtltNB6ZrU1TFmm9LAN2OZoVoczD83JraGcAkD2BabVprjUForCXE5kWb
/sTP6My9KZn1J/hPnuEbpPau63J/w1u28dWJLz4X/onSevUxnaPsXWc5f1K3iGqTTNbMNOUVA9xV
e9ASWXLkDiRVC6QcsnJkR1TlZgJzGLxduAjw93kDb5xincsKP+nvOdH6NkIelftL509tWRU4QDKF
aN36j8KcBOovx6Lp/p5YiPbIXp/BB6kjsfw2HfBxdcp0TF7lHloR47Kjd/sCyWbk7ugtWLN3Pccl
Bmciu/ORQzr+yK9ZQvhmMIjRI4BXhcdULWlEQQTUj7xLnwJYp6U6SgYJH1OCHP090n0z+r8Arj3v
0K19LK1TVfOYyrnxcyVHY+kZIRYk7sXHqyCbR2RmJstt6rp6WajaFb4CiE/oDe9kMxHRHqDZp25t
ChvG4H8YdRF6rIbyWx9xQPHqgH04Sm4QYpnb4+/cvJxyr7Qy3VhKgHPyzVF4jAMD5bPx5GXPTHSq
hsR4PnirTXlvgBUao93+qVw36bLy9W10pQ2EnTnEzaHGX51pfFaoZ1vKiWhc3v5LbkSByKzrEWq7
uTRtricDACLG80MngZA9UoV8iUbiHFq2HZClcZRAbtTET/Hj7agBwNQvsWj9jpRuvE8Yn0lb2RPR
qekT1c5gO9agCuHXZO08ByhCDZky78RLVW5c2mml5+GR7TWLtkNh1/jv0I6tXrfZCtn46BCnhhfq
sHA7NUuIQc8up0baxmYAXdWyozKF8CAyERwx2kJDMkOynRnvrdtZVQ/aaPKdEEkOy5O1BjuPLyls
FMS7LtBSTuQWYff54bhHqQrWpTMdhKiYTCqguQJ3ATt+VzaVDz059BKb/pnBpj5Ikd8sA3KZxynT
E/fTDEkYFzAD3pRm2gotbZCgYJwJwKrsMhe+N2AJhuA5Et13TRpB93JNlwBEu08NIlYJ1FTZEAFc
mDxvaRZjfb1iEeYualvatCuMgHNjCMn7TzgD98K0TDFMtwS3b5SIais2fDxLWXXSpe8VfEhS3mkz
NfIY3uNcb8KurrPgJ+sxdLgcD8t0+myeDgzwNnXELmGa/vtO7ut/Ti60ZymWqX7S7yDZ/ljGiWw5
aYRE0eNEaFIoa/ooRjOlaaTjiTmcfxN2MDBVx/pWfR8dXSvsXd+IGh3+3aAGU/yYKTHw4omxCiXt
PwdsH+fu4hzjG/vr6MTlDNRKpX4ZwSMKtVIHgDJynoFU7hW80kie2LBZDUqulcbtz+BtKfBY2ZM6
NW2ryCU2HA+1QE5TLD1yB44liKKq+06IyBLZ6W5akzdWTgNJCxdslT/V3rtKqMgErOH9xnd+zXje
BjaVOBMK8lZVzz06zIrAucg+i7DPSW5Fw49OeDf7Sg9r8hPTNKCLjtdp8ybOHNFor16lpBOwifw7
qVO4VT0fsBNg/iqHwspSUs+Z3a/UeNcYTFYBi1uirtpNfsaLWtBe9mYVXO49W6s2EQ02wz1aqzlO
hb2jVqonYaHF8NTD0LOnLQ/JyMy4DRxxrY6t8Exrb54TfVctoFyGgo/XNbVuqCOuBXyRntL2aSIp
W1Ur5KdQ+jRyCqccrZpE8EJ+i9o5Hah6lRyvWXnAIchXqARg42uv9W/N/QsX6vw601kgiyyLGp7/
o+dCzyAbkgUNxuBFl2iOZTIfo8XL+NBw0D2oCgVK7HT8KfyR3Du+tL7lmIGHIcoZ0T+1h7UJfjxW
RnhgzW5bCsjHSOPYvB9wrMk/x2cBfa3P5+WgLDbqqzN+3B7yHsbDWtLIwRYuqc3mZe4MfhE6QIfQ
CsseQxWaPK64b9IHxRHWpRRawHhAJwmZqdnfafB8cq4ACwexfWUR9ge048CR+kh/BBo2OR+c9M2r
v9pcFxr93ZAMxFrghcLIp0naceDpO/2BnMSSfzcMWI1gMXb0Y2zPPP3ZSpVlpGhHZjHgTEvAuwY5
BtDp3B9Sa+gWUjzXrFwuj7cBUQ7Tx//ZnZnKDMfZ1e/Z+WLRvsXg8IJ/PZEcbteOK1p0vSKI4iQj
yTuly4rbwahPY73CWT7eSIVjNby5DQAij0xPyo8xlxAx7mpbebMA+UW6s5ksoC/p9DSm9diAbKH4
VwZt+RSulCDKSLvO3eqcLfbIN1kIHFR6eWvoS/Iid57XJePu9PY+NPya2GHUk/e2Gjeso8MpmVbq
d3H+hIPVTN185fElsLDJU/8BEWeetJtMBeIA/PPj87M/4A7IBzDraDuwMYAttMStpce+TAVklrac
pRYSb4mSak6ee732pPlMqbiBMgfmbncCnc05IP//5Hx96qLw0yCz9EvtDiBW8x1w22hBDDgIRvgm
f6bB1h4s1UghBgG+g8X5PVN/3zAodDHs32NeQQJjVr7do/V40uJIwbnlgUepaQOar9xtUmuFvfBy
OVaeWCjq/n8p3s2O5JT2vddBXB5Q9IeVeVHfXN8Lvkk9Cu6LFsSUD+wR4PQxFtlQPHS1oHPs7VSu
6UG6TK8nZbg0caBLQVq1j3Vg6Uzme2PfnBICRg2KYfMf2Q4Iv56UF18DpQywaBCmpzrXQPN1dIsz
BkrJa4l9nxR9TzQ8bPVtGldOGTwqG8eqC6Uz5tuZTuQTTxjKXkZ7dMrNZ6LW9WVZwVEoIETmfpxC
JENAL5qyPLyqPgJJAcytgR+OsmowL7FRD5U2NcOaeZkInjpw5bxpa7n6M6adFbPks7zVGFOkV8mB
c0yjJ6rvgOHjql5R1bMp5UC4oMC/uWTSVcu20i4zNyqzI6UivB5mSoJFaGsdGya4Gn8oiV7hD5Tl
lgawtmlO0jo51am6tAFsQ6UA/suu9e+OiQDNB9QmYB/Y0aZaXDTTJaILPySLI45k9KZPfns+7AJr
DWE1wyU0saHJVVWRcRYh5nhNMiIlK5QtTOqbXa6/CR4f/OO0c4xfqVNvhSmc0o8+M1P3Rj2HRhhs
4yADBimNwA6Fs3h5o3EqNfpnIJygDlLhhYnrSIttX6EG2hCGwcchiTA0rW8cPGub/1DB4ZWppSai
pxs7UgcFQlEhNtcZHC7ol1Pnq/ZjS3dpIMhTi2P4EfNXpth/h8Kr9/fAv4rU9OJxV1IuT6F0Gd8Q
ZIdpC7j1bgNCFJ+I1AD4aj0gfQ0FHcWHrugoRtELlGct3SbW01+GYqtBmEhFMvULsMWFBFmym6d9
2XILIp8zIID0KhT1UrSGhVwRKxOQuKZ9xXkPU5S09saBiTEBwYp/auZ0nTjH6k7YAdblko/btvMw
/SmOI5xmn8GusC8xhoMCj7Mseeq8ACb5N0XpgOfDA9CxGJioeOIWt8+Hglfb+4wLw4YgHB6Uo5C+
s6QTbB8TioyghyJJGgGZxHtg0pv16JtYEhqxKuQgYHr142IET9ADXI6b5CNKoMD9fzM/TapqyIXe
tB3CGzLfiYo+7s7kT00LYHJiSwJ7RWvZcaSMOINB9VOiTiTph1l25IvTnPqMcXzCMIACwD50h6G3
/I+VBNuYJ0OlLUFffPwjuSrhfJw2MMGREfO2ADam3iXJOwrdka3orlBMfCrFIc40N9Quql3EhALR
HndCFDWVMWVxOhwBvNQmr/rX8Yc14of8N3/EbHqJYOm19i+EmEsVUvcsrBHqT63MJfg211gOU1bM
HVfgSmF3+mZMZ7E/wsx/Jrapkux2c1MtbEt1eLsQOhHW7xCLBpiyRLrWhPs8Rj8nGpJsYG8utnDR
Bmwzx/KCfQMLn/BqtMf49VvdjQnp8fbU2LIzfhS9R3t+w0cIfry1Kh+kKWCAZclUocI9IKrc3XxN
gITVQZsfDyjJ6gigLWqSMqwoPcRyc9Qoig+/B2SoroedYUCVU5DFbymx8v/Kcs7WYfomJh9JF8yg
GoN7k8TvbBVzEFaAij8OH7ktd1c+Enx7SzosELkpKeJ7gu6cdimJvhRuCLvVUznMyuOP0lJ9lgVB
xZL/VC5PSbnEgsmCoKJFTKhFTJJkVXjLnerlhKmiFPAyEeQYdEvq2ykHSYQzTD5RljGdes5xkC2Q
0nS+ctkj+FX63uZMjxcQnxhHgAsn3MQ1VFcLtjOzQdKoT/kF1rmyL7YZn//xhVIOwOs8mpJKbdUl
zuHIMe2Tj+bX+tLM86ZvIsJbRZzoCODm8xv21XZdSeKJ6RHdIaWKeVkkS3q8eqL+nYbXefEgxZDc
+1jOnt08QG/bYXZ1POSbjSRMGzjuWJBQSk4k3ijGM51/YqqfUZ33I4h1adpAQlh6NHB9YmnYa2xS
ffo95Tol73HM5SpzG+Nwailhfz9/NfUZYT1sLkF0BXNIy5de1K613flaIzWq6SQxWh0L++2TuQDV
kKUisOg/ppBNvSojBAsPGjPw2blD+GydUTC0lb5OvflC+hLjrZ4jpmMk6VUH2B/e/71EgnpHmxwC
9yt5LUJJ6iKyIL4k7hjKDCqZWS/KIRnd5Tfzz9n+RmM+do6kjCKEWUrwM8mG65LuonF/NY+nr3Di
S42vTW61sQGa+2rqBl1Brejw3m/RqgbiZPiv4rcN3dO05RZ10kQzvpab70br+mtO0hexvFv3Rrc6
Oh8ZbQF2A/w7iRzBM2ydc4LNsq9KCjQWJhyI1Tu2k2SYkIo7CbVm4+zJ5+CigRh8EoTnq+1Vihzi
/Eo+vvdCFpRELC/ct4ooawjko69s/ovJAOROEmHn6ydZr+7UAUZlfcHXUgfKgaTHgXgcjW5F9Vp6
HWP7ldo0juGa+R1HJftP69a14MsJA3aiLy3G0rlEjWRRPJFdfc6vDZcKUT74QLPGY3GTvEn7Ub47
RnH+JMS+uPWX9StIZElxExmxOB2eYfV3huLEhRX97naA16SgBQ1qJVJTj4r9CS7xMUgZ2IT87G5B
YPxI1qq1w730HEE32iUy2xoPWgKLPtSrI/mMnyjAaclyx701xiEj3WyPa0ajX+nPiJSKrQWs9BiO
B9vxW3bA83IZ4ZAKzZGLdyCmMlD/TLfnKjZ3FY0LyEvL28Rld9lDJprGE0pxvZzId3gJ0v8h1w4M
MABGc9WbGYVuoQHHm896z68D11nN5xFoD6t1Eln2QjShrwFyFnZeVVXS7ft1tWu9So678SJLf15g
7mEcsVyZ3JhBy49nlIx+K5fDH2WUvw8jxMaXEaL/0dUOYqwn5TcGHMBcf9ME4LkNN+2r46J2L308
PsIEjqR/7qncvWn3TxsyJ+xU8uUiqKdDcHTWJU+qBhCWlw6PX+K8ZdYDceULfjR1aAo2U/KjzKhy
+PFZh99r/PV/YQvsgKTEWI6h+qA1cXEf93B6qYDWmp2HdGQgoMRU/QdUI1iz75gEAmNgnIezBEY2
DFzFEO3+Bd7BCWv3tnPKnjrDrHM6d2w21yNbVKrauc4ZslAlKhTIOuBGq6SbUDdln4PJ05QV/SZ3
qijmBk+pAGjjEcYlce8cmNNPICJf9rL5RORu2szcbY2/zfHL5ouc99xbTx2AWgjRbN+etE4a8LVu
2YoK9y1n4HYi/8EsN1xzXyk/hvNMudZc9DHh+s9E4IURsS0dHzlGa9vlVQzdLbICYdwePAMM3MrN
JzVxHclotTGkKYF3HZ8vZNwCPgtC8UAUduMK7oiMVAGfGjzrLcOzRMinkwtHk2EfFOhga6jLMioI
WdhNTrtUPg+59NqNtk5/WEUTz2rbnGP8a9l5S2FbyDGtKPaGrZsY+qMyg+2xDOkychz3IaFCsis1
180aXnqA5GRR19LbgyuahSMfKnjnl9NDaxHlx0KQ6A5r65+oaZHcQ2mYODi5SLz3rU/oEHHdM/eD
uBojAyJIUQXhVHdmcm8erqV2IMFaTdSrMGYLl9T5QdfCLafUEI9cP0ijzjClCC+3JSVYli2NgypT
5YkpsBs4vlv+4G7rD77Kn7h8KhRbF/NTWBwicm24r2CLEib0CUnLeSZxROS7GeR7S6PjCUKiFsgC
vdf0CRteE8pjzZtI14npN8r08QIM/roqhRog/lXDVWKNz/+oYmLeatT/T1HdAtIRKWu7shKPsJb3
Cgj5s6THy01oZSVCVh0Em0HJ3lm5uiun1Ebv5MtLeVi2TtHw3uiII54qhC1d/juxMpissWo7urMv
Ryp5yLPGiEMkIzdrXxOUmC7ZeuJ7x/YryhDIfaKhB9zvdPy0w5TSnORLWveHzCf5eqzDJE7giC/o
FvNJUQO6AIpIypdmxPqwUemwL8cT8bcdUBZvbbFjCTpO2Z/GU3SvB9L3/g8b2nx11L4zZpNq9sww
XBvYgOXsVo94ZSh3s3Qw2XgFyb7U+ghz8ta3RkvDUOs8s/tfrQgbX1CsuqGL+lhf4e2ZasY7fAIT
8NagwAVTtw7u8AXBpbs/qa64pHtRlvgyKjCJbRzwDgGRb/Nk0/wQTM6ljB4xo1UVh4shjUKHIdxc
RKhGDFqVJ5iixLpuvpp2GHfBqkXZU2acmRgl19WdXSy2xFveG3jzf8j4Ce/Oj5kkgIDBNDcrU6F3
W85qKMCbaqGglqniLJkBxDLmqouIDCu/vjI8/wz29NSz0tVUpzmP0q7gVikMt3Pg+qQKCioKnj6o
4TtImjkzsPRJdRD+AdVzO1ggMAcM2bp/At2uNZrJ4pU770kiPs+ry+OwjAJylsTW8LLOGHeveh85
wBRbqiEvyHy/mHpHWEBFqIM6hpjEdHSNvIR/EqW170HQrTMrXtisySoqsepagVcpcMLvZ0QFsCyh
UCO103yyFSTlb9CytxqumWyNWHzNGaRcBzYlWlrfNOgOqBr5Nfzx8/sco6dfKtXJLtx0VjRIJ2VB
cKEAtXZG7Eu34NIE3zSI9cDmt2Cm24xqMGcIHg8DJW68q+aqKNX+dKByUcNPUevcEVlXFW1hgcQZ
X7pgNdwvaMR3gURbm43kqv5ZyKoVL8VHOFy01aH/j62Axs+DEJZ2ic3Ysu0/bevizKY28cqsmgEO
6Y2MCtJmCXslgc+mN5mL6mHl4GBqM4kVQ6aWoStGM0YBLCBPnHDDE4un2U4NsCpAmwYwkdX61ZQn
hLeffndfXfooRs+WFFDX3BY86jUS/mINrufS+bo6Mb/nbPvEBfs3VV2mTV6Nd7cS2HkrkQFIAYtZ
Wb2H6B5ZHrtjO1Lwa5vsZ0eJE9L9Iz2SOEVSpkZgeP2jX4VEx0ZyUzlM2t83Qm1YjziWjVMnX4CB
cRTL6oT/7e5HFlA0I1bmq9URD+xE641hoS6xbcUp+ZZnl0UMo0gJrQZr29HWdJPddKVamgauUjuM
QBfR3LuDHAwJFIjtX/QmmOjPH1LKKPzmaLEL/KgVywcGS+izxqEOFkBnWX6P/WK1t8hb3EeanqxL
qGghtWsdslA08hq2PQGBuEvK/0p1TxfOzceGGTdbBKoJhFtC8FR+thjESquDU+1sr6ZCsYOAfeaF
yzSptF1ygX2eGwDra1glQ8akwa6jM2WnRVgaEvoUnN3ieQrgKh802cbNDGSSOdIUakLK53vavGvK
ZSFZkPgbzLMbhBwTi5hdVgneuLG+prRmpRo6+lyf2vNI1Yhrtck2aI34fX5gjhq2W+MFAb52LZpv
duFl7VmsG/4Sjqc/gKHoRTFrHugA9fVerkHZuaGMyMAqe5zN/1xIZi3YV03xR75IeqCGR36VJEcA
aBgL3vOc9qoBubsr3A1BLK3tXwY8TWhU/45WTKC3maCsjlBS4AbnIq1meuVNdd9svsWmL27gQqf0
h97FZu8uzmpFMMWjfbaCzveb2S1N025HqF/q4dqbrnDxLfyvxX5WXM3k0Ux68raSCGRJa7+VBdzi
bLXDSu24r/m4Vv89/7Y2qkVlXaUMYoLcLd6Oaai1uUXSsCf+4rU1K0H+SZftn3BBlaG0XnQb9H/p
SVN589a6/nfxAh/NaiMHn2ZBCU518H7ANXyq9RzZCwr8HmQpFfFA2n5MbB8aRsg6h7bP53PZ5VYr
8RnCuMmNkMfN9nl/XQiDzRHVaAK2Fgibt2oph7fFDxqK3/QNIgLrT2kSTeSMh3zOy8W/6oUH1RYJ
Ux42E3M6zkUaQnyx/LEwsVgWRfmyNHuntYWTPdgHwgdAiCmEEOLmJbYX/X/+PWBAVa9jWldLo3Iq
vEFVqUQ5BjGD12LuqUTTaKT3WW6ruonkQ2AELMfQXE39jDc3z3YzY9Zxs/BhfnL3B5iGlbOCp1a6
ZQiR0DGJVLnci7YO7e/NJjrPSyPpd0bt3/tktFQIxEilBdO90UJrDGBQvO0HiNV3sXaJvTUzRKvz
eSsoedtPm+cEH3TD6IW3TeIvT4PGuJFWD+CZnA5IHNLL+hqZwoNyXn/7/a+WtlK+CMXknlaxPIaa
hd405DZhBqLuLVhIkMrtWHfUfgAj7F09SstBBeMHU3WZc71LSp15y/pgzjQipwE0FODl0Q1LZmgE
sWE/k9N9i/NlnRWLKWVgSy/craIn7wOAzHSNRlBl6jFqFlATc+2etPsxgCxidEvR3XntM1W7QC9H
MQVjdmqiS9ouqvBrxsD3Ivro/Mst2xxW3FLcPQ2z1itvqJe0bf+aY0g5yZw3gg6K034OUHoIIme8
Z8QWxvBVR0SSgA3PgRFJVYXDR8PWdFhOy4FN1VWgYndcS5QEnd5+blMw4VQ2ojFcxY9EjjYeJ8P3
MCOH8S7nrj9tu31vWFi1YsczFCnFKq7tbIlcJtPkH/+UB7VTUBr740B0lSFFsDhhv/CrBXN7FRrR
kMW5C4io6j0Wop7fHvqF2ne/IU4FOVBHF0aeEBzTBF/fG0metqpIboRX833P0Q3+JTtTJrmCJEQT
Z8Nm0uftlmxxKPNJtD+3YspyyMFnDTcZkoAfdjDfD6sMJ+IeJlBE4A+5mppTIH771Su+IOiXip9t
Apf0NOaTl4oTZYHvnm0UkJX+eI0VoS5QUTR91KicqB4lXC9mag8TooBqKyrrB0tOikoLzs8SBabS
XniLt/3PTbwNfIQVUYlaJjmzC6eFnpKMgqfZ3IGy313KwSvY5XoyhVbGaqp57zYo4W6BoBZrr6eu
B7Qem7z3pqFonRUdSZEYaREzVviFw6pjemeShGKpY89OHei/bsa7GLTLLywE7j8vvPKkqgBtTfrS
oysx2xiI5hLF2w/UE1fVx1HEfzLFCx/xkZ7VuYcXH+vhAVLcTqlaqLHg8KL1pvmAxFycxM7ui7DA
Djm6BiEOHcluf0aofeCpofoUm5gTs08eGZ5I6SuTKcv55Sp9Mvx8TsSdBxGc82omZ19sR1jEz/k5
BK2BZZdSGoBT4PrAeeHNlgecZCKxzFtvNPu+jvF6cjoZZAIqEzpSHYKCDQkytzr05kbUY3TIzTlD
1ponH2cKxuTcB6ibZgwX430f3cjZt9aWQNJ68TQGunaoiSWRcGtq5H12E/iSfB5YPFi0GsVGhf4z
RF7Q+pfhU72M1AemQOcxmrCKu0kRL2U+xXa7YhVjsscIHV/n+dGncTdLfvDGk7Q7ZfZJ5bKwIZkt
3Ga+KLOrAeJhPSvJOoJU/mTCmmDI4kSw9jlAipnqeyEYuKcuw7VD0We54Zr0FSC01hU38i47fVtd
Pv97AkB+6Gnc9YZhHqj133FQDW5DDoybnAc1SHLMLRXzDJ38IJVWWknxjI+rWrZapnUizJpVhH2m
ITSV8MatGFYie3DWOc0NJfJmsIbGF2Bh2nGLMU4tgFgdnuawGX2jNN47uThpA7EFzIokaYOPqOR7
ygQWdmw7aBx4WgISfYb4j5lZ+db9aC+pWL6rAy2MK26azsnnhsiDbIOwCTVAT2vvQTthclLEKcQk
fheJGEHPTEFsTfH/O/NuHkaSUp4BmZxYl0SQlKy+B6oeBF+4hHnPf7C3PONKOrb6mC06E3qsS7BQ
IWdSEWqc4hDvaNz4FpBkPj6h00tlTGXCP5AFQuGNbCXvnXld/kRIC+EW79CwZur2owN0Aqf4MDc+
inUybYWuxtUwATmrmkiYp0RWAnQD4yZP5Hbpr/o47tsE2GALNfjzT8wsiOCeFgF7Qk30wccPeysz
ciqhM9DT5SObSN/5m97lFFJ98I9L5Ecwzj1pP+K80ZncS39eodKH5G79LjurFBU/T3Z21wo+kofY
OrDBPDtGU4QUlkU7YCFTQynRz01uZMAjZxHKTTHE4gEFu0l1fTmNI43QqW7VlA57rzrDBQpkWYbw
vXjvNYTMfHQIH2euWkOpUZsJ7jdq+WOnInmm2Vd+vrsos9KJnChyIUFVNuC/VV5dwQ3Qu/HItG45
dPw8ayvbMlkBjP/IbygXL7txRfoCQED012xZpNk6X9RdC6PsdeCCP20RDIyh4vyCZbWqdkdgGBdD
fDjBjw8PBl0YZh5i+lQ1Z7U0xXfXi8TXNP0gz7442/B14TFgt9QtaSPmZ9+1R5JsU0jhjSf3ZLQw
Y2zXBNV/h43NCLWFllDmn98vhHZdb4qqeItK+zKGxoSDZIYzh+kFRUYYA3SoY/gZ+WZsbBvfOtrC
OCPeCqh/KtDOfLyJAcR8wY/RKVio4riSve6aop3wX0hyOcjbYTjp3VLBAsjDwdyE8yYQhkTqKsre
B32X7lEbJfNmzalU3VKNy2COQ362sTq47EXgEmpkv0CdkXZxt5brxcMxV4zGJZzdP35KvRY2vb4k
mq60JyaySuwfKbzp4XG+8gZ5XrTne+XcuHlXH1MZVgZSQVkDr78EIa3zIJ0llXQcvYqYr3uZ0X1K
0a9ry8/jqtWLfsc6Mr6LS4ufPXQCGV3dp7nCsPMfI8tAPu97OmOYEmIHBBChJg/HerkchYITrgxp
FCnzH6rvukqC1TZb7SOxb5hzrM3FkLJU4q82+QDxImuiVijZHReooNRbFK/nmFrEeKfRlrhkorbh
tER4P3VDMAsUpC7b+xTUOmI2rFKZKCUFcp0fJnv6c++n5t02EdHWC7ozuG7aqWBwc4tyrjPSNKIE
h0SI3FmWnfhwQ3YlLZ7Wv8A8RtstqgZsQhYDRgJuuLPxj7NncvdyOK+4x7aUoSBw3twKSMTRfBMg
XyaAYcly32Ilp7F/hxwcfwlOi9Gds3S8eHRNFgvD+Io/E+IBRfdsnV6pmfS0LoiXv0eSeqjqZ1Cd
TOnxGIY096+qmPI9s3V5nwYS155u7EkRCq9WqY8J1Tjke5aLbNNe1dSo4/+FlQE6lc/dO7IJU5+u
5sNrKyuTk6LaSgl2LtaZdsfW9teLlN1Szs3PwvCjiq4GCi0iB4iTX4p0GtbZKMX4oh5WYLz7UIAG
Sm33hTyMGiPA6Av89WD6q/UHx7/u0c0TsWMJnrP9yB+9RL0GZEunPV2ySToeaDRVrkNe0ics2+b6
0TIzP8K4/LcD0HfzT3AaOei9BQCwi7i5E5qIXw47kFL5kVlyXTukVwJPnvgEU2hyIBO/xx4BhaTl
hvBb9p3VjLvncrubNKPt9mQDgw8/Hkd1Z7dURD1ya2t9YhGdcr7sBS/SpSCWBFxzTJMOdWZaFwG2
tXKBzIa513NHZx5M9PXDYjvlfcW/HRxjn2yF4WMTsJoLNC6zviCOi/GLnj96KJhAdjNM/ZYWBEk7
b8HrvcOKteB6UeWb/G7Re3Llk0BlJiCOT3yoLFVLkN4bHIEkFQTD3qY0VmQo0A+Dq/lsluUpcSyf
BNlcAFeqYjmhh+rUxZlkxt3G+uwNgzXsED5yxJc63jpE9OahO3Lrsf6Yr8ysQlz5EO/tyGFo5cNh
zk08U6h0r8HPYrFDJpiPQVLo2iru1VHsaQ665MtQHSVCQSGfcCumfSkV67Z4xmJL8C9wYw/JVh5l
+7VfeWidpNwBKEc0mpOeQcaOxvSSnoCHAv9GW003mD6oZlhDdW+hFtJgemBPM1NswvpoNpS/u7tr
DR4NYXgDyIaUmXfy754whi7nUQ6MbNJDGhv1NtpSYVmePFxBA7rS6x6Ay6nCldRXSkq2zYtAgo0b
q5Ykfc1Nm/AyrwRTJelfX1dbYmw4w73sFRwuAUzZmRcjVdBSVIgUNkoVw+i4aahH82VoHMDACtys
vKXM42AX0KHEKv8O5tkCMrFFhpN5Siu882P5W3rZcVO9sT73SL34kkFHiPzxesm1SwPEEP+KcUKK
FocQdGI+LSqPx6SJ+gBK46wow1fHKLsCz1HbiqpKS9Fu05YLB93G4gclciVinR5++njYF5lrn/Ne
r1h8zWT7ymTOwAXm9TivxDsPkKSHTpqZYTdtA0LiODQAKXe2qm0MzxrSb1DaZcvZ6/stOARQWLJE
kyxHlilb3YVhsf7hwbtMEN8kJpvPll0A5jkqq4iNoHLx3Xc1JN8OPTfXdRCR9yA0XXeJ0y5S0yk8
iSYa7orr+xCQPVn/qrn/zllJop7wfiivKQlRbEyRhiJh0Bx3XXp6+koYAvUsdIa46sSehWS13f4E
RKfwJKKkMrk9hRT8JRhsbmMTC+Xr6i0ExcHiCEbkuEgJwqewm6hRaV3MY3IqhH3OW8hYWa663JuO
nX3ROEB2hentnEjd0pT12jSCkn9jf8GYsPz2z05vqZps028RgdyMo6tNquQx0o59vPxknzcbj2AG
WEoIYrBfbba7p56x4j6+Pz0rCOcyeUHr8R1x+15/UapIG1rGMwJfQytpF9zrpCHYQ7e5qDH1AUST
avumbyu/1YgviMu6AT0I03wDBU0Rq2/ird+XerXVjH0StFAJfJvCB9xXYl1Xdx5Yaha1adLXGYIE
sgIekzLh0MTQ1TeWIs1r1FNwi/Dzy7ile+G7WxawXqJj6q4//g1PoMQQy8s9yrmHWPhv7srgxp/l
9etAIxJoLrxVuHxMDQzaJJjyr//EG0WA12TPKz0GZJ85WFFFgKAsIc82SSErsDhrzu4TiOaiHCNC
sEC5u0egigwsrHxjLubJvvuI9YIZhsKcIp5pzAu4jKhSiqH18ygJK/gzD4v2h1Ctt6IcH8EKxtD+
gT/wCBkDdJoZM28GY5iknRb8pph8wxEf0738KmgmSZQ9Cx1Ns1OY56BrgBwqR9bAumJnYzKXsAx7
damAfTfdBfccVwuru7iR9XY1cV3n1ujF1yWfULAjmLp70LTkNo2ED9mherDMlaL1/T3DCn4SRzzw
D8EdMl6VIFnGRoqkNApO/F72rkQfaGxPeBrHaH7U43DqGRKLjf0h+r5uGoQxbS0VzBBMv2+emTyS
ANGxBgQZ+VtQNrEMs5BD8jPuGp4xGsOCevYmdaFtNw789PJ4l6ewOLWGK0zS2P2dFuapMMSoJlxa
UBSAcdwgi+11TKfxXRoOlqoxyjJPYcMftUS/+VVHJlMs/VmkPwZ6TRVkiTe+wLQiwyh+1yoyteRj
eE+AkPPa7KhBcEWDMVIB4PWN1sw7BC0CY53IYvUWqDY082Acvd0YgUT20Tn1PF7olDjyiaSWKtM4
VGLhsSmgk3Ws2ogw701CyVeMRTuyXyJs77qnC0/0ZYE7XMk5iUu/tcfqOS3aoeuxNgAUSKHNjFRT
KE5p9vutywYSpU6tvTIN2ssy2ghSKzebsUMewol+NEwULpJWXFeRt+FjOzkU93MYclL6XJU/5zhN
D/2HI3x5xr8WGxiLZrb2WvfxmTahgyhKSg6wuS0f3VSnnMot35iojhquZI+bIE8AXSL3f+ir3POM
w+LD9INTp9Hz4evermPImKMXyL7RXaBOLDFijb3th5j0KV1Qv/PIVlP13dkEp0eUkcfpjZLUDcjH
wGEgdIX8kVFQm/QAHTKWLQUCcHnZj/FtlkV/3HMulJ9/v85+Lmfb/zT6J9G7xOv2jI7DDZW7uyyz
rOSLjp+tlYWXYS9FnRUyKDiLmUgpasDTuC7KCDrc4Ohrk0WAqtP3TrqS6v3T66917315lt9uq1mW
YaZSuO4LIVIdUYigM1zDPVgc3hAJBwMTH7vm5/ZWqjSAkBAc9p+fMeyQUwBDTWTdAG3oiuDaJBXW
SgDaXpwXueQYr5ifrL6y02XDPJ1RCXXrtRDutf+hF9MxcShNAc27Cbm8RzQ69odb/e/TtJmAQoKn
YpOsi3lIE7ej4ZcxLnLISCGIMTV9bN5o1i9byAKq7M2NKst18ax4ubSE1fGz3X9Ff4a2WT09jniT
wIJIOateIk4UJNYAb2q7CsBTrEWmkYyGUbkC3oAjePoT3lxHRuj93r94WGDiFwvgnoIM9OaFs3Rp
HbOHuElK2tuLyLhAfcl8c6O4KgYLxYjDuXiPJX70+YiTX2Gpbo6WvOO9/0RpYDr0dnrW4io8EAUa
66Nxo9+MLWI8HhICX1q7d06QB06bWH4RLZfM/9NkFxSVdqq5gvFFEJ2/mNxjz3pL6kLbc3aCOzDY
3YMovCwBG3DD7ZWcBTxxnaUL/lMNSnSFuG4cQ4W09jsDkTnXg+FW8nUiScQIrIwWonjyE0aoKPM7
R17eq5Xz88ALnRwdosf2XJ9Tqr4y8KNo/Nj50G0HLVFvpgDz/WG/CiJ3rGlsk94zX5cox8Kpjb+O
u81kTyFwX3VF8n5JjZUmytFa/VZljvztTGqBlKJSRK2V6aHfbBDVDfgGyorY0qxtP6x10HI5zqQT
dY0TjiOJfPv3pq+Gsyy7NFJNgKuVvYH8a26L8nygRUPVXKx1zdxenZXIcM8Y8gEyFSUW5ArAfhbu
khX6cnrfPFK/1uLLdHHq5PO07SewlkUIGE6DCQZdw9Ue8oWhmHIkdMgUF27qiVMGA8BdoGMnFH9q
orTH1M3y8ucm3ii5PYGBmGGnLfeVZ4hE3KEYVGKHGbYwVlHTZXCkBz3G/Nt0YtiJHvdfZXDVoIvy
6AcQU7VJIt9IWB6LnxRgt1956HJcnPBvlqWgvChh4bwdktTY6kLxJKWV0w7Ae0QsKK6105C9Xv0v
xWi0R/8PE3thrIBUs/7fRyJe1hgMHD/Z0EVGl9UgXCcdaoq7JOOn5AXc0m7E1FEbBYW1tY2ftOZm
jB0z1NoOGxfllqH7r+WIoKq+n4VJ2r5rDVs4jNSAOvTEN0D4qe5J9X9nHnZwwo2cM00QONCR7DM0
FRoT0ICc5eBpjCu0xBN6yVJCYQZY8cmSayy30sIG1z3O5DHhy6QkgRZz8CKqdY3zJSkBP0jKzbB6
52wDtX74/zeT4XyEsJ0wiGvR2swuYItkthEHMIj9zrpnA3vZanxjW62XrQGOlC1nEo1Umw9eEYgq
zxxZQMh3X7leHafHWgA6gA7cFmdcspkdMEo5Gq6IQTZVE7KzOrEmWAFj2/CLaGvVay7c+Kfjl56P
xqsS6rVX7zbGJgs0bv12UnlzqylZZuSWOEIxF2HPB0OwMiHKxrYZCn6051C7z+a0vg81nd/ubB56
y8S/WqWhqB9En7bth7DZ4uN911iZ1ZLgFBo+44YZTiet/ELA2Ya14qQ7xkppJhNJMSzo2wnpDbdT
tj11wB2RZMZzkB+1lzUH1/gGFmVyGq6txA1iSHbJhqFTbYjAZJF+g9KDM1R1x5Mz7cLpdXHY+LeW
JdMp4nkinvfbUcknEE60FitO08PvYr13jYkOSq2DvhUzZCNJg+7ECgqiFlwO8Sn5gcnUKY+LP4dN
HvlaXnUUmMddju0m+9JaJJqYDbib89dIhffCSoX7HlhfdNoiqNggaEzqLVB/+WRP31gj18NTlLMI
ABBreL6ybDecwA69cethIkFplZPILQwA/GaRUwN79Ru1euCNbpgNYfbVAg1sRLJG/fs7+RiUKAlA
JhC7PsnsTv8IHXDSX7YT+SUnSlauIRV8uy0bxoYoCJTrpJ9c2M7+Sv1QznGEUOcmjW+zZZtDgQAk
GPsllRyVINnSDiVmtblMFCrNWUIqDeEbbhlRI+AIb2ppomANTGpDhFkXt5sJ4kX33SofPHj+0pkO
UozQuJLUdIiaj9GbpncZrePHdi0jbDRvDKEIS2RUiFmmG8JTdHRtEPXm4XL7BtiRli6SXBf14T5q
t2/mIQk7dEjwtiQcvpg8SYinygSs8INZVbwb1iuJoqKrGnJaenoW1yWr3flNs2P3oyYV8MZZdual
Ne0Xhl60FAd/g663sySAhJpcTpX/FwUiW9TZZDiezNqNnmxZR07bcyssRwc7JAWKAj8Er2v6zshW
uZ0+XiQ+eVxaoPuNO+tS4Lhx7G8z23YfW5JRtiN82ohcNMgZULYXvLu7hqKxf0NX4EMX7v42e3WT
qpySHx9Pmysy4XZni81ZQuR1GLRISmsAaC8syp9TlRD8HvXq6IokfxN3cUTC6Po4zEd8LExtn4TI
NNWLnFSit4Zsr9DOON8vdKuNP7+Z29uKdig/4l2gg4wYQ+pe0GTKb2BU0v/vZ9qZnBMWBnKDD3ki
tz8ETf0s/1HwPqQKzxZr5a+U5nC5IZ17qjcPaJn80ybZWhexRks98nANDuseI6MQ7DugTsYjfpWg
1TBOpmTD4OlmEe3uuxSs4g99zgry1ppGxtmZmeUFMT1TbUXIVJ1roUbs0MZpbNGTqWWQi6e0qhT3
Ge4P09202tKtMMlchXIyuVnosa99Rjsm359yxhuClOPAHgNy3wPMMQKEUrmU4uAByeqFEb0CEZT9
hqY2o3Qib5d3ft42JQrWttLSr2zKLUUqe4somw0Vr3DUjW14aQ6b0SkKk/NMYpHX+HsT5g/uK4T2
ya9oUNOUF/9dthF8tSx8gGT26mu7B8ed+B9Htjt75gwOWUlazDBTqssno3J+YsqDBHAcWHSHfNTs
yx59Wm6+T6pJwAm04L5KlLC9u0G7UY0L6/RNBsVAV+gUZaWLqU97b0iP0wNHF3ADLHzgyJqPbYsc
ND7yWlHgOcgGecSu6Grlvng7mdl+iPZUbpzDT39ivygANcd6Z1julMrlcDbLUv/GWaLetMj14gFP
F9zg2eLtmkMD9+ELV5zTnH3yX3Dlc/yKKk8EMhGYgbFDHgXCUMH6IcfMp3tONT8P4W6ciyUCQj4j
M/zHC8Tv6TS72ZObPSVWgbxmObxpWDU8iT1s3Nwk7KS4ONIes1YKsjRXb3Nukm/NcVui7+CXW579
mactWDOF/gGIi9+efkqQaETesTUK4fSoZjjTvpjhNmRvsL6STgPslchI0zj7LeWPgowXHgTNOWxk
f2/p0SlCtGSHj9Eei4jF47vfqn0W19/eXafujrTVqAnuGTF9/qWz2dRKzmkbI6yRoGDOqg9M/o2d
ioLtX4hPvOpINe/Ghnl5owOf+jNVo2md2hcP3IQ6QAXNsD40rwn62uS2nESttgm9LGqJ/tEXOY1l
UbiJJfvfpEAc3Wz7+/VVhZyo71RHQRyA24u5ZUcJZU3xn0RYFMb2bIXizM9Q+DotvALsFTcT1sxo
l+AiqmVVEvjc1fxhoGG1SqO5AmC0U9P55m/86OWUHrn7n2L9QG/7xxyXt7KBM6JwF8wQVe6VDjTI
5SoKyWeG5TTeyyXMYOTUVe7RY71XoTAdukoD29JJR+37khcy/JML8OAaf9mXUjbHRYoDDYqY5hlF
CtpmLPfXeu6nKotZgiJ2xO3Qo2+evVNbcZ9tYjyT7NyixRzP7rEaEQkq0kmPEjregCh8rPOwc+tK
pliynxA/iDhF1OHjQSsK+zVRpNV7xfWCHsSCaqBz5+wc09lNxJfYYIC4gRPU2ZfZpUekuAnjNGOj
Uxm0Lu+lTZZ1GKIrfSADzfd08sXqldRd+2GlD5/Pxw+7IT5fLTY9RWLoa9vntVPa3BtnLfcMt1Jy
o3TbOOjlAUjZisvysXSfqA6NQq6RNfXM9+2gnzHNju9nJeRBNbNm+4vcalgQGaKE+2dNnAlqOVLr
3oL9UnpTYasH+zWcsfIxRMUu4J7a3ZhzK+sv9nE7zG8ZNHMCJY5G6folPbhZCh7GelxVs/7zJS3I
WpzmRhbQmJkSzhvvFxofczp4CxUDlUs1vkIvmYpEdnXJrKQUEZFk1oAIijt+5SKBJkBBlRmsLb75
Pqgk36M9Wyei9d4ldsSDRcKsPEIqI6e3k0BaCkCRMi/FNY4nn3nu3GE01JP98zgTv2Ag8+9DOOvG
Hd86pBYoKbcFv07kmtGW7tCk9kcAkq8DKfo000E9KjV+BC+P2cbHF2+BSWqfJEJWtnP3fZl755BI
IibH5pDuEGUJvgWsWVrlbVtDvChBnVT5aO6R+B6gMuz1u4eJS8szMh/rCceOKpJhb+YMBhYNLqHZ
Em0VONeEen73dgtSGhSGGq8Sq9LatlNY6Fy2er3bPwtu/qZH67jOWrK+/bPWiprXmnTH0oQ42cyp
7LYsy1YE7G6boA250ud/fSUCEQ33vLKVMMGSkoyOx8K849RGv36mI9tRVrsdmyEnDKAFcw4Ic56F
Wa9fyeLBw3yTNehP4WL10fCvSXOEW7Al+5fN/XzJOlfdDtoEFBr9fA541ehKjdzHBvAYUqslivO0
d2b5FQA5fufyWOGN40KcZjCyZQmC8IZa5bl6qzQFEDAOrUj8aODRxqBrF+4fGa0oFTzDf7vjBQvl
+W46q+b7Bpqu+HkBpKnGI2PepY1jTMyk4X0RXveVAd99IDx6uwNyiW57KFt2g1iHp/YIIMh6QX4y
sJhJUW7vxqCwJjn7opCko7BmEkkR3CHYHUZu+p5Fj8tap/pmMvMJRqvUwBI5tRlzfDOgH2AirZbU
QVwS8lBm7VlcpJEaqlrA410vMOXcDHiLuvHiVdpWFRWFngvaL14ywm2NEuk+h5hsV5v3MgPKAKOy
kPrmI7Chg47OjYY+6i5uy3DgOvw8lKWyKYusLxJ+U+n9P96UO3NHw4tbODFzFsEckHLF4SNre9HJ
EfOeswQdiHRCnZV0xR2BnxscXqSIicrIhqTXoxeUGFXD6G87J1X0E85AbU0uYzWhIMQlAIMKYzBQ
WKLoqrXFcXQt+W5DMk3wIK3ovr5Gfa/gCshZH9Giswrcg7jQ5Zvd8+m6pXW+pWsIzBoiaD9aQQDX
ehJoUqJwdt60gbKLPyobP6e2D0kLHC9D5iEwy1Hs21ycbNHc8dyJDBJweussT8Q5iUv4uCBkGExP
uChrczoDLFd5m2JvLhOfRN3p2nCw19j2vSnhtt9/8XZCDq4nQom4FxG65drVP6u5mcPjEcxeUfWt
e95DfhC5hyaQ4nNNv//jkEGaX2njTjERAr+gK5woHglERMQTlvRmhNy/49jdaZiHk30RdoSP/MtI
J81t2EWYn+9r2wieYRKNK7XahuHZrisS6Uvt7d1KffGvefKhq7W/0J1Zht+5gqaN1KCLwX1KhHAn
89YjAi07ml63HXq9Y0gFfNEX4/JLWbEZ3MpjT6Vgj5zJ7XRXzgdgwjGIny+KYuPPgjOkoeA9DvYm
7SEL7aSjbwq0yiqD0PkTNGCHLIiCBiY4qeETp0to6pKEy7RRU4AuFDfLfqfAcJNhaV5mx9MbUiqD
gASz/CLFpHUkGv+xJ3COFTYH1jU3M2ScfXYTlQp9e6j9zY4E8PjpyC3t1AI99/i0fB3h/SAvpU7t
BWqo/gw4S3KclFLotEELyLFxkkBT4344P4yDHK9UIgB8x50hFopGxjS5YCon8r/6ul/YLFZlUysz
r+bhvpGGoL6ZkNubRnj8avCCRa5gVzcv5266DCHubA2z8OE8IzPyEbcL+LqO5ZYgdzVCvir9yPtA
u5pWbtyZMCdYEHXL/8rPMnqUBDPJ2z9iQCVmCugGrujhltBgorZkqfKS7DQ19NpJlYpEVUMv9EIB
VAECgqEZ7LhHJQSsV3Oz8XgnAx3RFNb75X6jz7W9Avbfen9zkwP0Psk6HwCXj4CEUAYaY/98cirf
9B7DzHYk5nQp5xnWMVImVuzTpAI8XRj4BSYv2YZewSVirBsDZz6nclgSROb2Ehzpr37fgGH/J+vN
hXnnD3uNJJnTKghdd/ZprDSf1FsaOkvOqfo0A4OOufnQyHj3BhLhMqCh5/Fea+hK9jdGoJ8ax8+p
p2f8wwr3InYt00AT3airWlesHjE9ErqfVqoWlgkFBBApWOurUZW6oK0WMpucKpg9KdyHukBDiCPy
qX0PN4xr95+9VLrY6yYqiYJMcyI6ENFZQ8Y5SDEMsnezdU/WRGl3ZeXui0CHswpcPr097p9nRQqa
/6hyRUZ/cYIFq8nDCAM7KiFkvFUJbkFDZEGScuzr7AstZkqE2VE+iI+eLQTYs+tg2dARBz8YWhV6
m+MET1qsm89MCAedsA3pit0LzxfymubBvVFYQiCfzXjBvxGafttTtTQL4hzOwwLEOVIThnyJldef
ZjPwHovJU2Hrx+VZR25R4FSK6lWKZ+vumFL3vG3N+qw9dbvy/pIskIRGt+/GvVAWxxiiJYf5Xuf/
77tYbN4p2QmmtaMn8+5Wkafpj22lIe0yjkPYvOKgFTzuUGQMya2Vm+GfKIWuAIv82WuAJ1FxOH1/
4IN/zCJs8S0qzQDOJgYY/LqkPPRm1MWRQBNbFqNLynog63cozuj6d24j5v5dfB33fjIJ6FenDPWR
bPCIB5Bm3ZWBicNKZRGlyO5EHXKKD7ERdNk1lsspVY172C6LGFItCuvqLmGixyx49hddjhCq/cjo
Mk/lkrXlGLsaQernaV8Z0Q9tqu9ISc3aallB2gE2Os0l367adEWLwtuVnkqja8ljFgbNMMjbQIzy
jVI7rUoReiKYf5vpwQqT5yGqU2VqPHReySzYSqaWdCn4uMCmsbpnjCdwOKoKHdxYG0pJZpju5mGr
GPznwdkWHU8pkRvkE7U0vuYEmoRdUSBXdtqb9UOCMrAqhF9YNoF3Vi/ug1tWVnga8O4vq7OdyWLg
W4vLgEX2VogegnXD8W4H1MCY0p7Z1gqaK+xMyPt5wbLq5sNFOafZcicakNCldaFbC4J2kVwGjvJ3
9opRY8cgshNOcKFcLrmdCZJH2t+wry8P+xL6EERVqjE3nPWwdy9RrZxuQPdCX7odB7V+kBfUP/mn
ORnSVA/jGnkrg5ZUcwKPgFCh2y+xHraXml8QRQnwUP/5MHtUvmVKFK6B/WMT+OvTV8+YcDGP0Eoy
pP8qunZwUCDRc9VphIrUnKMkj4FfRcEryGKyqIR+CIbL9koFP6LUSKRrXlbY4JwVkFHx+rbCAP6R
lQOT0iHW7jYzsLT9DVvXdh9wHN5I6WwLxjRlFKskeVDXOkKXByNAihRwObVVL7wSodcFBXzZ96NZ
3VEGwWl841/hYT7aXuc7dL+QUb0xfjTBpwuKVku3y+S2r9iDr50hLkOSBRgfGigB3hYwbQyXSQ6V
GKm+a8Ae80mzR9CydjemHd6DTLp9rb5h9qKkZ09zhx8qvmz6Kko0SmmN1Gyra6mTsODMl9VRfd+R
dsuxGQ1baoDhIVB4SsoEViKXT1XL02/uii9x/ZKaIrSCRmi708HuVue0tos4ur0w4D3vcEYG4dMx
4ALTLV54TAQxOAK4Xex09DhWDRCpD3wlNDLt99iePo8GhthABh5bqGZe9We4gUrcu5LJ58P3o6fU
mbaFYW+3ZvbngurpgDWJ1fXIsK/LwtYjzC8aPOIZ5YqKXYscT8QlGJ1HsB3Y3JzeTYqDwOmdGLjn
LlNPzaNtRWxJ6OmMRMC83Q5VRI4Y+DnAWJgUQ1QLlC/KYclMrglR7sbhDsR2t/8r82y289LKT1DA
8yeYwU6C3MrvN7rEIFxRkYwKWGsVwxGlIP1OL0XuOxDgXAq9c7J6aXaSPFhltco9/VWjhQtPdbF5
v4w5qqkYRjRVcOPJe57LBZNPsjc6mBrb7RM6a+7m7sqiyI5KFHezKIVfh2D+Z3YgTYrswfDbhXnd
mRjq9Vg+rUasOnhSsq+9+auEy6s7xSKCIJgRdTJNBwCMw3wZx2hi8pDRCNtiDQP+YBpbzCdmAuzW
nfJvd7FgVrnJBv3Pt03lYMG+CZGPWFG0I1pGHPGRtaXsM5FFrbezKhAj1OdQ8T3LPnS841fLngUc
+ftlMTEuXsrLNg9avUVtqkjt2Z9qp4mwLkRjsEUJQZDu79JeurVBCvqr2QvC0bBmjBuOzRkNt28K
soXYxzSaSlx4sMwfxLo0HndylZv5fpOjyoVsvnUprc6mEffHAH6TK5HmUVMwawFXlTPnbgjcjyLD
Fz6ar9MWAnhVUnh/dBPymAirgEB9mcbR5BqcSeAv4v5gIRa3N7T761WzxFf1kvpDSg/qmb2/6GLC
cCh5pgJrk5Yt3QgE/CCEB8VwvOXvOFbI/kyvCSYmJwKQSVtqOwcuCOxWXgJIPGuX1A8rfkiUSMD2
k9Mof2ZtvfzUglNG2kUsGayrIYY0XSfAn/GyvidH+Rg36Cfmmy4CrJc0mkF7XRLz4wXjmNHlZkFd
C3+v7/EY+3H6DdvdjmPcTA8UDyecuh3U+w3oJNfY/6d9JBoXuSo1/gLbnoLNuV8xEMpJEKuJvPFs
BHKyTbzwWB1Ty+kRlKuYwwurZDqAy/n+Z+Yp80QClui0dGlJWa3IPC3QjaLIPw1KNZZCmEGsSo91
rB7/O5e7pSA1KZLMayXLbIjy5LPvI8h1Rs0x2+7WUs2nNehqqGIsZq/hLs4SivfSqzUdcy04we/9
1ARp22N/O0REWlN7QOJUfe43dgjSnLkU43ShnFmLG8G6b0jRTYMjzVL4F9uX2xAPLwZDtkT5CpKZ
R2l8VN3nUnzL9fGdmJf6UdeLIRb+S81KzJbJCislkJqXsZ4oCNwMq26FVElKNqR4m0QewTZRkoY3
xkaT4d1aSAztmKIe0LWRZvjNsZBRTP59p/pDtCZyazsJEGbJxx3g/nsV6Jop3DEV4Df9s0w2rV5h
Ke1ZCZJEUbOIqqmoVAxrn78j6GjrfmI7rIf8+W76fBwdDfJDzvW9bQj03yIWVw5RdgFPJHxk8suq
sneu8hZjy0JcohtRhnGZb3YdjEhVvN5x+qOWnfyUIuWJmNdk48Kmujea9c41b/+wvYlN1vs/xcwB
iOtzB6CcJX029DE6ZcGHi2HmEE9V7XZQfnxXNV12SdQPPm5H1+MoqFQiUZrZjvm4CyVxpGVwLS9s
ieAYRhVw2T/smyt1LR7bqtLoNvN/qSUnNP+l8K5iMAVJCboLoQxR6R33zG6bx756AkOD2GyRPzg5
z8FFYFaGNXsTb3pxp0Vt8njsoW0xuoA+5bB11TXGU6EP2LyomQjzajuUbUQKU85AfX+xR9INCdg7
bCMGt0Ubw//ERka0m2SFTa8QeoJHc6YfF4nLO4sJNDM3nxAftsyqsuLTFtCJjvztqHjNZo6N7/5E
FCVLqwvzhwAHbEFBK7QKd5WDkcYRSh0CR+CXDWaFHxHTEmUQBDszIgDOFc8NBackGNpPRXRYiTOS
zk0FI4qgstxGMkaN2hDSetQnN4cam2ewEdhSYG71Xo+D7PbEBWAfraMPtlmOE17qfkgWM05i0Ama
c7MiPZXo92cVZczMSZRMwKbx39lClceaHVUfnnTzoJQ6VrPTxtClw23u2zhDBLQdCgB90D3QbBEU
aa5/MNxqyqMLWptb12KGVYk/irhAeajfK0kBphA04fpNklvEMl4l4Vtf62XSe3/3WPXZrNk1D/kq
71Zor4zVLO4guN6t23/7Dc532pAYslzHctezwIj61+JMDDiVoVGREqKoy64SEfcOZBvoX1/6g8gJ
0QdMtqZ6h2ZC02iUveWPDcff7X5g0A3j82rOXvs4eq62bWsK2QCfAZd2eOECevcIacuq5ZjCO/ja
dG3uQ7zXEh2kEDzRjsONmN3xjh3ZU9hBccGbofMQgnSD9LOO58CvDnHg23DRFHT5VioNVmOqoYXM
zeoCssX+gEv5LjnFR6t9suXwdmTkKqqoIyoSqu1peVSr1A2QKirqccIE6l3FO89DAB8Arihyr0hg
6W1cSaG5klJeAl4AeKLXbCSdVlTFfcs3quJQzavBdxLOG+cwNcUPWkTH9Te9rB8QoqzvKb/Dc774
OfObpD1EDcaUzs+KSOUgxhxuZ/VJ8Du5WWCStLOd+dlxQRSzme7C/s4+4a27XgkRLABv6lUnCtXV
6S/RkWb/LpGUkRQZpXGm2tc2HQDPcJRonCWI5xAbWyttWpCOaP4YyDAVY5Z3ux7Rp386WDz8ExT4
xwsMRLn4Lhexaypl2kSmTX3eCCUpaSKg3EhtYWiSzGCr9SXMc1gg6LfXxN9zqe/X9w2ujo66bzGD
kEySO4qq62oFLrzht7rP+MuiDDax+SejGjIsMkq1yhvdVBtrFsFXLmxl0HZnWyc8lUhPqMJ5TeEQ
gntgt1tqKWEbDGvVX2UAgjVOBRcC7MaGyEzR4wyU6Q6YIZBCpkNK8hFaLs3FngZ5Z/QonwSeQ//h
ecsJCTxMVUEPpYRBha3shKaMQveAz1Hqz2hbpffiXeW0wRBAAUk8fPRyTesUTLzed6vSFR4f/5qf
5em1iSD4EfhRu/4c27Tt0XU4q+mxzQDrXgLdJde86xauoK+Sdr5F62fjN4mFG8zgLJygo2Dl0D4H
+1yrKRL8HOhMMg==
`protect end_protected
